
module sin
(
    input [9:0] theta,     //10 bits of precision, first 3 are integer part
    output [15:0] out
);

parameter [0:9][15:0] ROM = {
16'b0000000000000000,
16'b0000000001111111,
16'b0000000011111111,
16'b0000000101111111,
16'b0000000111111111,
16'b0000001001111111,
16'b0000001011111111,
16'b0000001101111111,
16'b0000001111111111,
16'b0000010001111111,
16'b0000010011111110,
16'b0000010101111110,
16'b0000010111111101,
16'b0000011001111101,
16'b0000011011111100,
16'b0000011101111011,
16'b0000011111111010,
16'b0000100001111001,
16'b0000100011111000,
16'b0000100101110111,
16'b0000100111110101,
16'b0000101001110011,
16'b0000101011110010,
16'b0000101101110000,
16'b0000101111101110,
16'b0000110001101011,
16'b0000110011101001,
16'b0000110101100110,
16'b0000110111100011,
16'b0000111001100000,
16'b0000111011011100,
16'b0000111101011001,
16'b0000111111010101,
16'b0001000001010001,
16'b0001000011001101,
16'b0001000101001000,
16'b0001000111000011,
16'b0001001000111110,
16'b0001001010111000,
16'b0001001100110011,
16'b0001001110101101,
16'b0001010000100110,
16'b0001010010100000,
16'b0001010100011001,
16'b0001010110010001,
16'b0001011000001010,
16'b0001011010000010,
16'b0001011011111001,
16'b0001011101110001,
16'b0001011111100111,
16'b0001100001011110,
16'b0001100011010100,
16'b0001100101001010,
16'b0001100110111111,
16'b0001101000110100,
16'b0001101010101001,
16'b0001101100011101,
16'b0001101110010001,
16'b0001110000000100,
16'b0001110001110111,
16'b0001110011101001,
16'b0001110101011011,
16'b0001110111001101,
16'b0001111000111110,
16'b0001111010101110,
16'b0001111100011110,
16'b0001111110001110,
16'b0001111111111101,
16'b0010000001101100,
16'b0010000011011010,
16'b0010000101001000,
16'b0010000110110101,
16'b0010001000100001,
16'b0010001010001101,
16'b0010001011111001,
16'b0010001101100100,
16'b0010001111001110,
16'b0010010000111000,
16'b0010010010100001,
16'b0010010100001010,
16'b0010010101110010,
16'b0010010111011001,
16'b0010011001000000,
16'b0010011010100110,
16'b0010011100001100,
16'b0010011101110001,
16'b0010011111010110,
16'b0010100000111010,
16'b0010100010011101,
16'b0010100100000000,
16'b0010100101100001,
16'b0010100111000011,
16'b0010101000100011,
16'b0010101010000011,
16'b0010101011100011,
16'b0010101101000001,
16'b0010101110011111,
16'b0010101111111101,
16'b0010110001011001,
16'b0010110010110101,
16'b0010110100010001,
16'b0010110101101011,
16'b0010110111000101,
16'b0010111000011110,
16'b0010111001110110,
16'b0010111011001110,
16'b0010111100100101,
16'b0010111101111011,
16'b0010111111010001,
16'b0011000000100101,
16'b0011000001111001,
16'b0011000011001101,
16'b0011000100011111,
16'b0011000101110001,
16'b0011000111000001,
16'b0011001000010010,
16'b0011001001100001,
16'b0011001010101111,
16'b0011001011111101,
16'b0011001101001010,
16'b0011001110010110,
16'b0011001111100010,
16'b0011010000101100,
16'b0011010001110110,
16'b0011010010111111,
16'b0011010100000111,
16'b0011010101001110,
16'b0011010110010101,
16'b0011010111011010,
16'b0011011000011111,
16'b0011011001100011,
16'b0011011010100110,
16'b0011011011101000,
16'b0011011100101001,
16'b0011011101101010,
16'b0011011110101001,
16'b0011011111101000,
16'b0011100000100110,
16'b0011100001100011,
16'b0011100010011111,
16'b0011100011011010,
16'b0011100100010101,
16'b0011100101001110,
16'b0011100110000111,
16'b0011100110111110,
16'b0011100111110101,
16'b0011101000101011,
16'b0011101001100000,
16'b0011101010010100,
16'b0011101011000111,
16'b0011101011111001,
16'b0011101100101010,
16'b0011101101011011,
16'b0011101110001010,
16'b0011101110111001,
16'b0011101111100110,
16'b0011110000010011,
16'b0011110000111110,
16'b0011110001101001,
16'b0011110010010011,
16'b0011110010111100,
16'b0011110011100100,
16'b0011110100001010,
16'b0011110100110000,
16'b0011110101010101,
16'b0011110101111010,
16'b0011110110011101,
16'b0011110110111111,
16'b0011110111100000,
16'b0011111000000000,
16'b0011111000011111,
16'b0011111000111110,
16'b0011111001011011,
16'b0011111001110111,
16'b0011111010010011,
16'b0011111010101101,
16'b0011111011000110,
16'b0011111011011111,
16'b0011111011110110,
16'b0011111100001101,
16'b0011111100100010,
16'b0011111100110111,
16'b0011111101001010,
16'b0011111101011101,
16'b0011111101101110,
16'b0011111101111111,
16'b0011111110001110,
16'b0011111110011101,
16'b0011111110101010,
16'b0011111110110111,
16'b0011111111000010,
16'b0011111111001101,
16'b0011111111010110,
16'b0011111111011111,
16'b0011111111100111,
16'b0011111111101101,
16'b0011111111110011,
16'b0011111111110111,
16'b0011111111111011,
16'b0011111111111101,
16'b0011111111111111,
16'b0011111111111111,
16'b0011111111111111,
16'b0011111111111110,
16'b0011111111111011,
16'b0011111111111000,
16'b0011111111110011,
16'b0011111111101110,
16'b0011111111100111,
16'b0011111111100000,
16'b0011111111011000,
16'b0011111111001110,
16'b0011111111000100,
16'b0011111110111000,
16'b0011111110101100,
16'b0011111110011110,
16'b0011111110010000,
16'b0011111110000001,
16'b0011111101110000,
16'b0011111101011111,
16'b0011111101001101,
16'b0011111100111001,
16'b0011111100100101,
16'b0011111100001111,
16'b0011111011111001,
16'b0011111011100010,
16'b0011111011001010,
16'b0011111010110000,
16'b0011111010010110,
16'b0011111001111011,
16'b0011111001011111,
16'b0011111001000001,
16'b0011111000100011,
16'b0011111000000100,
16'b0011110111100100,
16'b0011110111000011,
16'b0011110110100001,
16'b0011110101111110,
16'b0011110101011010,
16'b0011110100110101,
16'b0011110100001111,
16'b0011110011101000,
16'b0011110011000001,
16'b0011110010011000,
16'b0011110001101110,
16'b0011110001000100,
16'b0011110000011000,
16'b0011101111101100,
16'b0011101110111110,
16'b0011101110010000,
16'b0011101101100001,
16'b0011101100110000,
16'b0011101011111111,
16'b0011101011001101,
16'b0011101010011010,
16'b0011101001100110,
16'b0011101000110001,
16'b0011100111111100,
16'b0011100111000101,
16'b0011100110001110,
16'b0011100101010101,
16'b0011100100011100,
16'b0011100011100010,
16'b0011100010100110,
16'b0011100001101010,
16'b0011100000101110,
16'b0011011111110000,
16'b0011011110110001,
16'b0011011101110010,
16'b0011011100110001,
16'b0011011011110000,
16'b0011011010101110,
16'b0011011001101011,
16'b0011011000100111,
16'b0011010111100011,
16'b0011010110011101,
16'b0011010101010111,
16'b0011010100010000,
16'b0011010011001000,
16'b0011010001111111,
16'b0011010000110101,
16'b0011001111101011,
16'b0011001110100000,
16'b0011001101010100,
16'b0011001100000111,
16'b0011001010111001,
16'b0011001001101011,
16'b0011001000011011,
16'b0011000111001011,
16'b0011000101111011,
16'b0011000100101001,
16'b0011000011010111,
16'b0011000010000100,
16'b0011000000110000,
16'b0010111111011011,
16'b0010111110000110,
16'b0010111100110000,
16'b0010111011011001,
16'b0010111010000001,
16'b0010111000101001,
16'b0010110111010000,
16'b0010110101110110,
16'b0010110100011100,
16'b0010110011000001,
16'b0010110001100101,
16'b0010110000001000,
16'b0010101110101011,
16'b0010101101001101,
16'b0010101011101111,
16'b0010101010001111,
16'b0010101000101111,
16'b0010100111001111,
16'b0010100101101110,
16'b0010100100001100,
16'b0010100010101001,
16'b0010100001000110,
16'b0010011111100010,
16'b0010011101111110,
16'b0010011100011001,
16'b0010011010110011,
16'b0010011001001101,
16'b0010010111100110,
16'b0010010101111111,
16'b0010010100010111,
16'b0010010010101110,
16'b0010010001000101,
16'b0010001111011011,
16'b0010001101110001,
16'b0010001100000110,
16'b0010001010011010,
16'b0010001000101111,
16'b0010000111000010,
16'b0010000101010101,
16'b0010000011101000,
16'b0010000001111001,
16'b0010000000001011,
16'b0001111110011100,
16'b0001111100101100,
16'b0001111010111100,
16'b0001111001001100,
16'b0001110111011011,
16'b0001110101101001,
16'b0001110011110111,
16'b0001110010000101,
16'b0001110000010010,
16'b0001101110011111,
16'b0001101100101011,
16'b0001101010110111,
16'b0001101001000011,
16'b0001100111001110,
16'b0001100101011000,
16'b0001100011100011,
16'b0001100001101101,
16'b0001011111110110,
16'b0001011101111111,
16'b0001011100001000,
16'b0001011010010000,
16'b0001011000011000,
16'b0001010110100000,
16'b0001010100101000,
16'b0001010010101111,
16'b0001010000110101,
16'b0001001110111100,
16'b0001001101000010,
16'b0001001011001000,
16'b0001001001001101,
16'b0001000111010010,
16'b0001000101010111,
16'b0001000011011100,
16'b0001000001100000,
16'b0000111111100100,
16'b0000111101101000,
16'b0000111011101100,
16'b0000111001101111,
16'b0000110111110010,
16'b0000110101110101,
16'b0000110011111000,
16'b0000110001111011,
16'b0000101111111101,
16'b0000101101111111,
16'b0000101100000001,
16'b0000101010000011,
16'b0000101000000101,
16'b0000100110000110,
16'b0000100100001000,
16'b0000100010001001,
16'b0000100000001010,
16'b0000011110001011,
16'b0000011100001100,
16'b0000011010001100,
16'b0000011000001101,
16'b0000010110001110,
16'b0000010100001110,
16'b0000010010001110,
16'b0000010000001111,
16'b0000001110001111,
16'b0000001100001111,
16'b0000001010001111,
16'b0000001000001111,
16'b0000000110001111,
16'b0000000100001111,
16'b0000000010001111,
16'b0000000000001111,
16'b1111111110001111,
16'b1111111100001111,
16'b1111111010001111,
16'b1111111000001111,
16'b1111110110010000,
16'b1111110100010000,
16'b1111110010010000,
16'b1111110000010000,
16'b1111101110010000,
16'b1111101100010001,
16'b1111101010010001,
16'b1111101000010010,
16'b1111100110010010,
16'b1111100100010011,
16'b1111100010010100,
16'b1111100000010101,
16'b1111011110010110,
16'b1111011100010111,
16'b1111011010011000,
16'b1111011000011010,
16'b1111010110011011,
16'b1111010100011101,
16'b1111010010011111,
16'b1111010000100001,
16'b1111001110100011,
16'b1111001100100110,
16'b1111001010101001,
16'b1111001000101011,
16'b1111000110101111,
16'b1111000100110010,
16'b1111000010110110,
16'b1111000000111001,
16'b1110111110111101,
16'b1110111101000010,
16'b1110111011000110,
16'b1110111001001011,
16'b1110110111010000,
16'b1110110101010110,
16'b1110110011011100,
16'b1110110001100010,
16'b1110101111101000,
16'b1110101101101110,
16'b1110101011110101,
16'b1110101001111101,
16'b1110101000000100,
16'b1110100110001100,
16'b1110100100010101,
16'b1110100010011101,
16'b1110100000100110,
16'b1110011110110000,
16'b1110011100111001,
16'b1110011011000100,
16'b1110011001001110,
16'b1110010111011001,
16'b1110010101100101,
16'b1110010011110000,
16'b1110010001111101,
16'b1110010000001001,
16'b1110001110010110,
16'b1110001100100100,
16'b1110001010110010,
16'b1110001001000000,
16'b1110000111001111,
16'b1110000101011111,
16'b1110000011101110,
16'b1110000001111111,
16'b1110000000010000,
16'b1101111110100001,
16'b1101111100110011,
16'b1101111011000101,
16'b1101111001011000,
16'b1101110111101011,
16'b1101110101111111,
16'b1101110100010100,
16'b1101110010101001,
16'b1101110000111110,
16'b1101101111010100,
16'b1101101101101011,
16'b1101101100000010,
16'b1101101010011010,
16'b1101101000110011,
16'b1101100111001100,
16'b1101100101100101,
16'b1101100011111111,
16'b1101100010011010,
16'b1101100000110110,
16'b1101011111010010,
16'b1101011101101110,
16'b1101011100001100,
16'b1101011010101010,
16'b1101011001001000,
16'b1101010111100111,
16'b1101010110000111,
16'b1101010100101000,
16'b1101010011001001,
16'b1101010001101011,
16'b1101010000001110,
16'b1101001110110001,
16'b1101001101010101,
16'b1101001011111010,
16'b1101001010011111,
16'b1101001001000101,
16'b1101000111101100,
16'b1101000110010011,
16'b1101000100111100,
16'b1101000011100101,
16'b1101000010001110,
16'b1101000000111001,
16'b1100111111100100,
16'b1100111110010000,
16'b1100111100111101,
16'b1100111011101010,
16'b1100111010011000,
16'b1100111001000111,
16'b1100110111110111,
16'b1100110110101000,
16'b1100110101011001,
16'b1100110100001011,
16'b1100110010111110,
16'b1100110001110010,
16'b1100110000100111,
16'b1100101111011100,
16'b1100101110010010,
16'b1100101101001001,
16'b1100101100000001,
16'b1100101010111010,
16'b1100101001110011,
16'b1100101000101101,
16'b1100100111101001,
16'b1100100110100101,
16'b1100100101100001,
16'b1100100100011111,
16'b1100100011011110,
16'b1100100010011101,
16'b1100100001011101,
16'b1100100000011111,
16'b1100011111100001,
16'b1100011110100100,
16'b1100011101100111,
16'b1100011100101100,
16'b1100011011110010,
16'b1100011010111000,
16'b1100011001111111,
16'b1100011001001000,
16'b1100011000010001,
16'b1100010111011011,
16'b1100010110100110,
16'b1100010101110010,
16'b1100010100111110,
16'b1100010100001100,
16'b1100010011011011,
16'b1100010010101010,
16'b1100010001111011,
16'b1100010001001100,
16'b1100010000011111,
16'b1100001111110010,
16'b1100001111000110,
16'b1100001110011011,
16'b1100001101110001,
16'b1100001101001000,
16'b1100001100100000,
16'b1100001011111001,
16'b1100001011010011,
16'b1100001010101110,
16'b1100001010001010,
16'b1100001001100111,
16'b1100001001000100,
16'b1100001000100011,
16'b1100001000000011,
16'b1100000111100011,
16'b1100000111000101,
16'b1100000110101000,
16'b1100000110001011,
16'b1100000101110000,
16'b1100000101010101,
16'b1100000100111100,
16'b1100000100100011,
16'b1100000100001100,
16'b1100000011110101,
16'b1100000011011111,
16'b1100000011001011,
16'b1100000010110111,
16'b1100000010100101,
16'b1100000010010011,
16'b1100000010000010,
16'b1100000001110011,
16'b1100000001100100,
16'b1100000001010110,
16'b1100000001001010,
16'b1100000000111110,
16'b1100000000110011,
16'b1100000000101010,
16'b1100000000100001,
16'b1100000000011001,
16'b1100000000010011,
16'b1100000000001101,
16'b1100000000001000,
16'b1100000000000101,
16'b1100000000000010,
16'b1100000000000000,
16'b1100000000000000,
16'b1100000000000000,
16'b1100000000000001,
16'b1100000000000011,
16'b1100000000000111,
16'b1100000000001011,
16'b1100000000010000,
16'b1100000000010111,
16'b1100000000011110,
16'b1100000000100110,
16'b1100000000110000,
16'b1100000000111010,
16'b1100000001000101,
16'b1100000001010010,
16'b1100000001011111,
16'b1100000001101101,
16'b1100000001111100,
16'b1100000010001101,
16'b1100000010011110,
16'b1100000010110000,
16'b1100000011000011,
16'b1100000011011000,
16'b1100000011101101,
16'b1100000100000011,
16'b1100000100011010,
16'b1100000100110010,
16'b1100000101001100,
16'b1100000101100110,
16'b1100000110000001,
16'b1100000110011101,
16'b1100000110111010,
16'b1100000111011000,
16'b1100000111110111,
16'b1100001000010111,
16'b1100001000111000,
16'b1100001001011010,
16'b1100001001111101,
16'b1100001010100000,
16'b1100001011000101,
16'b1100001011101011,
16'b1100001100010010,
16'b1100001100111001,
16'b1100001101100010,
16'b1100001110001100,
16'b1100001110110110,
16'b1100001111100001,
16'b1100010000001110,
16'b1100010000111011,
16'b1100010001101001,
16'b1100010010011001,
16'b1100010011001001,
16'b1100010011111010,
16'b1100010100101100,
16'b1100010101011110,
16'b1100010110010010,
16'b1100010111000111,
16'b1100010111111101,
16'b1100011000110011,
16'b1100011001101011,
16'b1100011010100011,
16'b1100011011011100,
16'b1100011100010110,
16'b1100011101010001,
16'b1100011110001101,
16'b1100011111001010,
16'b1100100000000111,
16'b1100100001000110,
16'b1100100010000101,
16'b1100100011000110,
16'b1100100100000111,
16'b1100100101001001,
16'b1100100110001100,
16'b1100100111001111,
16'b1100101000010100,
16'b1100101001011001,
16'b1100101010011111,
16'b1100101011100110,
16'b1100101100101110,
16'b1100101101110111,
16'b1100101111000000,
16'b1100110000001011,
16'b1100110001010110,
16'b1100110010100010,
16'b1100110011101111,
16'b1100110100111100,
16'b1100110110001011,
16'b1100110111011010,
16'b1100111000101010,
16'b1100111001111010,
16'b1100111011001100,
16'b1100111100011110,
16'b1100111101110001,
16'b1100111111000101,
16'b1101000000011001,
16'b1101000001101111,
16'b1101000011000101,
16'b1101000100011011,
16'b1101000101110011,
16'b1101000111001011,
16'b1101001000100100,
16'b1101001001111110,
16'b1101001011011000,
16'b1101001100110011,
16'b1101001110001111,
16'b1101001111101011,
16'b1101010001001000,
16'b1101010010100110,
16'b1101010100000101,
16'b1101010101100100,
16'b1101010111000100,
16'b1101011000100100,
16'b1101011010000101,
16'b1101011011100111,
16'b1101011101001010,
16'b1101011110101101,
16'b1101100000010000,
16'b1101100001110101,
16'b1101100011011010,
16'b1101100100111111,
16'b1101100110100101,
16'b1101101000001100,
16'b1101101001110100,
16'b1101101011011100,
16'b1101101101000100,
16'b1101101110101101,
16'b1101110000010111,
16'b1101110010000001,
16'b1101110011101100,
16'b1101110101010111,
16'b1101110111000011,
16'b1101111000101111,
16'b1101111010011100,
16'b1101111100001010,
16'b1101111101111000,
16'b1101111111100110,
16'b1110000001010101,
16'b1110000011000101,
16'b1110000100110101,
16'b1110000110100101,
16'b1110001000010110,
16'b1110001010001000,
16'b1110001011111001,
16'b1110001101101100,
16'b1110001111011110,
16'b1110010001010010,
16'b1110010011000101,
16'b1110010100111001,
16'b1110010110101110,
16'b1110011000100011,
16'b1110011010011000,
16'b1110011100001110,
16'b1110011110000100,
16'b1110011111111010,
16'b1110100001110001,
16'b1110100011101000,
16'b1110100101100000,
16'b1110100111011000,
16'b1110101001010000,
16'b1110101011001001,
16'b1110101101000001,
16'b1110101110111011,
16'b1110110000110100,
16'b1110110010101110,
16'b1110110100101000,
16'b1110110110100011,
16'b1110111000011110,
16'b1110111010011001,
16'b1110111100010100,
16'b1110111110001111,
16'b1111000000001011,
16'b1111000010000111,
16'b1111000100000100,
16'b1111000110000000,
16'b1111000111111101,
16'b1111001001111010,
16'b1111001011110111,
16'b1111001101110101,
16'b1111001111110010,
16'b1111010001110000,
16'b1111010011101110,
16'b1111010101101100,
16'b1111010111101011,
16'b1111011001101001,
16'b1111011011101000,
16'b1111011101100110,
16'b1111011111100101,
16'b1111100001100100,
16'b1111100011100100,
16'b1111100101100011,
16'b1111100111100010,
16'b1111101001100010,
16'b1111101011100001,
16'b1111101101100001,
16'b1111101111100001,
16'b1111110001100000,
16'b1111110011100000,
16'b1111110101100000,
16'b1111110111100000,
16'b1111111001100000,
16'b1111111011100000,
16'b1111111101100000,
16'b1111111111100000
};

assign out = ROM[theta];

endmodule