
module cos
(
    input [9:0] theta,     //10 bits of precision, first 3 are integer part (unsigned)
    output [15:0] out      //16 bits of precision, first 2 are integer part (signed)
);

parameter ADDR_WIDTH = 10;
parameter DATA_WIDTH =  16;
logic [9:0] addr_reg;

parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
16'sb0100000000000000,
16'sb0011111111111111,
16'sb0011111111111110,
16'sb0011111111111011,
16'sb0011111111111000,
16'sb0011111111110011,
16'sb0011111111101110,
16'sb0011111111100111,
16'sb0011111111100000,
16'sb0011111111010111,
16'sb0011111111001110,
16'sb0011111111000011,
16'sb0011111110111000,
16'sb0011111110101011,
16'sb0011111110011110,
16'sb0011111110001111,
16'sb0011111110000000,
16'sb0011111101101111,
16'sb0011111101011110,
16'sb0011111101001011,
16'sb0011111100111000,
16'sb0011111100100011,
16'sb0011111100001110,
16'sb0011111011111000,
16'sb0011111011100000,
16'sb0011111011001000,
16'sb0011111010101111,
16'sb0011111010010100,
16'sb0011111001111001,
16'sb0011111001011101,
16'sb0011111001000000,
16'sb0011111000100001,
16'sb0011111000000010,
16'sb0011110111100010,
16'sb0011110111000001,
16'sb0011110110011111,
16'sb0011110101111100,
16'sb0011110101011000,
16'sb0011110100110011,
16'sb0011110100001101,
16'sb0011110011100110,
16'sb0011110010111110,
16'sb0011110010010101,
16'sb0011110001101100,
16'sb0011110001000001,
16'sb0011110000010101,
16'sb0011101111101001,
16'sb0011101110111011,
16'sb0011101110001101,
16'sb0011101101011110,
16'sb0011101100101101,
16'sb0011101011111100,
16'sb0011101011001010,
16'sb0011101010010111,
16'sb0011101001100011,
16'sb0011101000101110,
16'sb0011100111111000,
16'sb0011100111000010,
16'sb0011100110001010,
16'sb0011100101010010,
16'sb0011100100011000,
16'sb0011100011011110,
16'sb0011100010100011,
16'sb0011100001100111,
16'sb0011100000101010,
16'sb0011011111101100,
16'sb0011011110101101,
16'sb0011011101101110,
16'sb0011011100101101,
16'sb0011011011101100,
16'sb0011011010101010,
16'sb0011011001100111,
16'sb0011011000100011,
16'sb0011010111011110,
16'sb0011010110011001,
16'sb0011010101010011,
16'sb0011010100001011,
16'sb0011010011000011,
16'sb0011010001111010,
16'sb0011010000110001,
16'sb0011001111100110,
16'sb0011001110011011,
16'sb0011001101001111,
16'sb0011001100000010,
16'sb0011001010110100,
16'sb0011001001100110,
16'sb0011001000010111,
16'sb0011000111000110,
16'sb0011000101110110,
16'sb0011000100100100,
16'sb0011000011010010,
16'sb0011000001111110,
16'sb0011000000101011,
16'sb0010111111010110,
16'sb0010111110000001,
16'sb0010111100101010,
16'sb0010111011010011,
16'sb0010111001111100,
16'sb0010111000100100,
16'sb0010110111001010,
16'sb0010110101110001,
16'sb0010110100010110,
16'sb0010110010111011,
16'sb0010110001011111,
16'sb0010110000000011,
16'sb0010101110100101,
16'sb0010101101000111,
16'sb0010101011101001,
16'sb0010101010001001,
16'sb0010101000101001,
16'sb0010100111001001,
16'sb0010100101101000,
16'sb0010100100000110,
16'sb0010100010100011,
16'sb0010100001000000,
16'sb0010011111011100,
16'sb0010011101111000,
16'sb0010011100010010,
16'sb0010011010101101,
16'sb0010011001000111,
16'sb0010010111100000,
16'sb0010010101111000,
16'sb0010010100010000,
16'sb0010010010100111,
16'sb0010010000111110,
16'sb0010001111010100,
16'sb0010001101101010,
16'sb0010001011111111,
16'sb0010001010010100,
16'sb0010001000101000,
16'sb0010000110111011,
16'sb0010000101001110,
16'sb0010000011100001,
16'sb0010000001110011,
16'sb0010000000000100,
16'sb0001111110010101,
16'sb0001111100100101,
16'sb0001111010110101,
16'sb0001111001000101,
16'sb0001110111010100,
16'sb0001110101100010,
16'sb0001110011110000,
16'sb0001110001111110,
16'sb0001110000001011,
16'sb0001101110011000,
16'sb0001101100100100,
16'sb0001101010110000,
16'sb0001101000111100,
16'sb0001100111000111,
16'sb0001100101010001,
16'sb0001100011011011,
16'sb0001100001100101,
16'sb0001011111101111,
16'sb0001011101111000,
16'sb0001011100000001,
16'sb0001011010001001,
16'sb0001011000010001,
16'sb0001010110011001,
16'sb0001010100100000,
16'sb0001010010100111,
16'sb0001010000101110,
16'sb0001001110110100,
16'sb0001001100111010,
16'sb0001001011000000,
16'sb0001001001000101,
16'sb0001000111001011,
16'sb0001000101010000,
16'sb0001000011010100,
16'sb0001000001011001,
16'sb0000111111011101,
16'sb0000111101100001,
16'sb0000111011100100,
16'sb0000111001101000,
16'sb0000110111101011,
16'sb0000110101101110,
16'sb0000110011110000,
16'sb0000110001110011,
16'sb0000101111110101,
16'sb0000101101110111,
16'sb0000101011111001,
16'sb0000101001111011,
16'sb0000100111111101,
16'sb0000100101111110,
16'sb0000100100000000,
16'sb0000100010000001,
16'sb0000100000000010,
16'sb0000011110000011,
16'sb0000011100000100,
16'sb0000011010000101,
16'sb0000011000000101,
16'sb0000010110000110,
16'sb0000010100000110,
16'sb0000010010000110,
16'sb0000010000000111,
16'sb0000001110000111,
16'sb0000001100000111,
16'sb0000001010000111,
16'sb0000001000000111,
16'sb0000000110000111,
16'sb0000000100000111,
16'sb0000000010000111,
16'sb0000000000000111,
16'sb1111111110000111,
16'sb1111111100000111,
16'sb1111111010000111,
16'sb1111111000001000,
16'sb1111110110001000,
16'sb1111110100001000,
16'sb1111110010001000,
16'sb1111110000001000,
16'sb1111101110001000,
16'sb1111101100001001,
16'sb1111101010001001,
16'sb1111101000001010,
16'sb1111100110001010,
16'sb1111100100001011,
16'sb1111100010001100,
16'sb1111100000001101,
16'sb1111011110001110,
16'sb1111011100001111,
16'sb1111011010010000,
16'sb1111011000010010,
16'sb1111010110010011,
16'sb1111010100010101,
16'sb1111010010010111,
16'sb1111010000011001,
16'sb1111001110011100,
16'sb1111001100011110,
16'sb1111001010100001,
16'sb1111001000100100,
16'sb1111000110100111,
16'sb1111000100101010,
16'sb1111000010101110,
16'sb1111000000110010,
16'sb1110111110110110,
16'sb1110111100111010,
16'sb1110111010111111,
16'sb1110111001000100,
16'sb1110110111001001,
16'sb1110110101001110,
16'sb1110110011010100,
16'sb1110110001011010,
16'sb1110101111100000,
16'sb1110101101100111,
16'sb1110101011101110,
16'sb1110101001110101,
16'sb1110100111111101,
16'sb1110100110000101,
16'sb1110100100001101,
16'sb1110100010010110,
16'sb1110100000011111,
16'sb1110011110101000,
16'sb1110011100110010,
16'sb1110011010111100,
16'sb1110011001000111,
16'sb1110010111010010,
16'sb1110010101011101,
16'sb1110010011101001,
16'sb1110010001110101,
16'sb1110010000000010,
16'sb1110001110001111,
16'sb1110001100011101,
16'sb1110001010101011,
16'sb1110001000111001,
16'sb1110000111001000,
16'sb1110000101011000,
16'sb1110000011100111,
16'sb1110000001111000,
16'sb1110000000001001,
16'sb1101111110011010,
16'sb1101111100101100,
16'sb1101111010111110,
16'sb1101111001010001,
16'sb1101110111100101,
16'sb1101110101111001,
16'sb1101110100001101,
16'sb1101110010100010,
16'sb1101110000111000,
16'sb1101101111001110,
16'sb1101101101100101,
16'sb1101101011111100,
16'sb1101101010010100,
16'sb1101101000101100,
16'sb1101100111000101,
16'sb1101100101011111,
16'sb1101100011111001,
16'sb1101100010010100,
16'sb1101100000101111,
16'sb1101011111001100,
16'sb1101011101101000,
16'sb1101011100000110,
16'sb1101011010100100,
16'sb1101011001000010,
16'sb1101010111100010,
16'sb1101010110000001,
16'sb1101010100100010,
16'sb1101010011000011,
16'sb1101010001100101,
16'sb1101010000001000,
16'sb1101001110101011,
16'sb1101001101001111,
16'sb1101001011110100,
16'sb1101001010011001,
16'sb1101001001000000,
16'sb1101000111100110,
16'sb1101000110001110,
16'sb1101000100110110,
16'sb1101000011011111,
16'sb1101000010001001,
16'sb1101000000110100,
16'sb1100111111011111,
16'sb1100111110001011,
16'sb1100111100111000,
16'sb1100111011100101,
16'sb1100111010010011,
16'sb1100111001000011,
16'sb1100110111110010,
16'sb1100110110100011,
16'sb1100110101010100,
16'sb1100110100000111,
16'sb1100110010111010,
16'sb1100110001101101,
16'sb1100110000100010,
16'sb1100101111010111,
16'sb1100101110001110,
16'sb1100101101000101,
16'sb1100101011111101,
16'sb1100101010110101,
16'sb1100101001101111,
16'sb1100101000101001,
16'sb1100100111100100,
16'sb1100100110100000,
16'sb1100100101011101,
16'sb1100100100011011,
16'sb1100100011011010,
16'sb1100100010011001,
16'sb1100100001011001,
16'sb1100100000011011,
16'sb1100011111011101,
16'sb1100011110100000,
16'sb1100011101100100,
16'sb1100011100101000,
16'sb1100011011101110,
16'sb1100011010110100,
16'sb1100011001111100,
16'sb1100011001000100,
16'sb1100011000001101,
16'sb1100010111010111,
16'sb1100010110100011,
16'sb1100010101101110,
16'sb1100010100111011,
16'sb1100010100001001,
16'sb1100010011011000,
16'sb1100010010100111,
16'sb1100010001111000,
16'sb1100010001001001,
16'sb1100010000011100,
16'sb1100001111101111,
16'sb1100001111000011,
16'sb1100001110011001,
16'sb1100001101101111,
16'sb1100001101000110,
16'sb1100001100011110,
16'sb1100001011110111,
16'sb1100001011010001,
16'sb1100001010101100,
16'sb1100001010001000,
16'sb1100001001100100,
16'sb1100001001000010,
16'sb1100001000100001,
16'sb1100001000000001,
16'sb1100000111100001,
16'sb1100000111000011,
16'sb1100000110100110,
16'sb1100000110001001,
16'sb1100000101101110,
16'sb1100000101010100,
16'sb1100000100111010,
16'sb1100000100100010,
16'sb1100000100001010,
16'sb1100000011110100,
16'sb1100000011011110,
16'sb1100000011001010,
16'sb1100000010110110,
16'sb1100000010100011,
16'sb1100000010010010,
16'sb1100000010000001,
16'sb1100000001110010,
16'sb1100000001100011,
16'sb1100000001010110,
16'sb1100000001001001,
16'sb1100000000111101,
16'sb1100000000110011,
16'sb1100000000101001,
16'sb1100000000100000,
16'sb1100000000011001,
16'sb1100000000010010,
16'sb1100000000001101,
16'sb1100000000001000,
16'sb1100000000000100,
16'sb1100000000000010,
16'sb1100000000000000,
16'sb1100000000000000,
16'sb1100000000000000,
16'sb1100000000000001,
16'sb1100000000000100,
16'sb1100000000000111,
16'sb1100000000001011,
16'sb1100000000010001,
16'sb1100000000010111,
16'sb1100000000011111,
16'sb1100000000100111,
16'sb1100000000110000,
16'sb1100000000111011,
16'sb1100000001000110,
16'sb1100000001010010,
16'sb1100000001100000,
16'sb1100000001101110,
16'sb1100000001111101,
16'sb1100000010001110,
16'sb1100000010011111,
16'sb1100000010110001,
16'sb1100000011000101,
16'sb1100000011011001,
16'sb1100000011101110,
16'sb1100000100000100,
16'sb1100000100011100,
16'sb1100000100110100,
16'sb1100000101001101,
16'sb1100000101100111,
16'sb1100000110000011,
16'sb1100000110011111,
16'sb1100000110111100,
16'sb1100000111011010,
16'sb1100000111111001,
16'sb1100001000011001,
16'sb1100001000111010,
16'sb1100001001011100,
16'sb1100001001111111,
16'sb1100001010100011,
16'sb1100001011001000,
16'sb1100001011101101,
16'sb1100001100010100,
16'sb1100001100111100,
16'sb1100001101100101,
16'sb1100001110001110,
16'sb1100001110111001,
16'sb1100001111100100,
16'sb1100010000010001,
16'sb1100010000111110,
16'sb1100010001101100,
16'sb1100010010011011,
16'sb1100010011001100,
16'sb1100010011111101,
16'sb1100010100101111,
16'sb1100010101100010,
16'sb1100010110010110,
16'sb1100010111001010,
16'sb1100011000000000,
16'sb1100011000110111,
16'sb1100011001101110,
16'sb1100011010100110,
16'sb1100011011100000,
16'sb1100011100011010,
16'sb1100011101010101,
16'sb1100011110010001,
16'sb1100011111001110,
16'sb1100100000001011,
16'sb1100100001001010,
16'sb1100100010001001,
16'sb1100100011001010,
16'sb1100100100001011,
16'sb1100100101001101,
16'sb1100100110010000,
16'sb1100100111010011,
16'sb1100101000011000,
16'sb1100101001011101,
16'sb1100101010100100,
16'sb1100101011101011,
16'sb1100101100110011,
16'sb1100101101111011,
16'sb1100101111000101,
16'sb1100110000001111,
16'sb1100110001011011,
16'sb1100110010100111,
16'sb1100110011110011,
16'sb1100110101000001,
16'sb1100110110001111,
16'sb1100110111011111,
16'sb1100111000101111,
16'sb1100111001111111,
16'sb1100111011010001,
16'sb1100111100100011,
16'sb1100111101110110,
16'sb1100111111001010,
16'sb1101000000011111,
16'sb1101000001110100,
16'sb1101000011001010,
16'sb1101000100100001,
16'sb1101000101111000,
16'sb1101000111010000,
16'sb1101001000101001,
16'sb1101001010000011,
16'sb1101001011011110,
16'sb1101001100111001,
16'sb1101001110010100,
16'sb1101001111110001,
16'sb1101010001001110,
16'sb1101010010101100,
16'sb1101010100001011,
16'sb1101010101101010,
16'sb1101010111001010,
16'sb1101011000101010,
16'sb1101011010001011,
16'sb1101011011101101,
16'sb1101011101010000,
16'sb1101011110110011,
16'sb1101100000010111,
16'sb1101100001111011,
16'sb1101100011100000,
16'sb1101100101000110,
16'sb1101100110101100,
16'sb1101101000010011,
16'sb1101101001111010,
16'sb1101101011100010,
16'sb1101101101001011,
16'sb1101101110110100,
16'sb1101110000011101,
16'sb1101110010001000,
16'sb1101110011110010,
16'sb1101110101011110,
16'sb1101110111001010,
16'sb1101111000110110,
16'sb1101111010100011,
16'sb1101111100010001,
16'sb1101111101111111,
16'sb1101111111101101,
16'sb1110000001011100,
16'sb1110000011001100,
16'sb1110000100111100,
16'sb1110000110101100,
16'sb1110001000011101,
16'sb1110001010001111,
16'sb1110001100000000,
16'sb1110001101110011,
16'sb1110001111100110,
16'sb1110010001011001,
16'sb1110010011001100,
16'sb1110010101000001,
16'sb1110010110110101,
16'sb1110011000101010,
16'sb1110011010011111,
16'sb1110011100010101,
16'sb1110011110001011,
16'sb1110100000000010,
16'sb1110100001111000,
16'sb1110100011110000,
16'sb1110100101100111,
16'sb1110100111011111,
16'sb1110101001010111,
16'sb1110101011010000,
16'sb1110101101001001,
16'sb1110101111000010,
16'sb1110110000111100,
16'sb1110110010110110,
16'sb1110110100110000,
16'sb1110110110101010,
16'sb1110111000100101,
16'sb1110111010100000,
16'sb1110111100011100,
16'sb1110111110010111,
16'sb1111000000010011,
16'sb1111000010001111,
16'sb1111000100001011,
16'sb1111000110001000,
16'sb1111001000000101,
16'sb1111001010000010,
16'sb1111001011111111,
16'sb1111001101111100,
16'sb1111001111111010,
16'sb1111010001111000,
16'sb1111010011110110,
16'sb1111010101110100,
16'sb1111010111110010,
16'sb1111011001110001,
16'sb1111011011110000,
16'sb1111011101101110,
16'sb1111011111101101,
16'sb1111100001101100,
16'sb1111100011101011,
16'sb1111100101101011,
16'sb1111100111101010,
16'sb1111101001101010,
16'sb1111101011101001,
16'sb1111101101101001,
16'sb1111101111101000,
16'sb1111110001101000,
16'sb1111110011101000,
16'sb1111110101101000,
16'sb1111110111101000,
16'sb1111111001101000,
16'sb1111111011101000,
16'sb1111111101101000,
16'sb1111111111101000,
16'sb0000000001101000,
16'sb0000000011101000,
16'sb0000000101101000,
16'sb0000000111101000,
16'sb0000001001101000,
16'sb0000001011100111,
16'sb0000001101100111,
16'sb0000001111100111,
16'sb0000010001100111,
16'sb0000010011100110,
16'sb0000010101100110,
16'sb0000010111100110,
16'sb0000011001100101,
16'sb0000011011100100,
16'sb0000011101100011,
16'sb0000011111100011,
16'sb0000100001100010,
16'sb0000100011100000,
16'sb0000100101011111,
16'sb0000100111011110,
16'sb0000101001011100,
16'sb0000101011011010,
16'sb0000101101011000,
16'sb0000101111010110,
16'sb0000110001010100,
16'sb0000110011010001,
16'sb0000110101001111,
16'sb0000110111001100,
16'sb0000111001001001,
16'sb0000111011000101,
16'sb0000111101000010,
16'sb0000111110111110,
16'sb0001000000111010,
16'sb0001000010110110,
16'sb0001000100110001,
16'sb0001000110101100,
16'sb0001001000100111,
16'sb0001001010100010,
16'sb0001001100011100,
16'sb0001001110010110,
16'sb0001010000010000,
16'sb0001010010001001,
16'sb0001010100000010,
16'sb0001010101111011,
16'sb0001010111110011,
16'sb0001011001101011,
16'sb0001011011100011,
16'sb0001011101011010,
16'sb0001011111010001,
16'sb0001100001001000,
16'sb0001100010111110,
16'sb0001100100110100,
16'sb0001100110101010,
16'sb0001101000011111,
16'sb0001101010010011,
16'sb0001101100000111,
16'sb0001101101111011,
16'sb0001101111101111,
16'sb0001110001100010,
16'sb0001110011010100,
16'sb0001110101000110,
16'sb0001110110111000,
16'sb0001111000101001,
16'sb0001111010011010,
16'sb0001111100001010,
16'sb0001111101111001,
16'sb0001111111101001,
16'sb0010000001010111,
16'sb0010000011000110,
16'sb0010000100110011,
16'sb0010000110100000,
16'sb0010001000001101,
16'sb0010001001111001,
16'sb0010001011100101,
16'sb0010001101010000,
16'sb0010001110111010,
16'sb0010010000100100,
16'sb0010010010001101,
16'sb0010010011110110,
16'sb0010010101011110,
16'sb0010010111000110,
16'sb0010011000101101,
16'sb0010011010010100,
16'sb0010011011111001,
16'sb0010011101011111,
16'sb0010011111000011,
16'sb0010100000100111,
16'sb0010100010001011,
16'sb0010100011101101,
16'sb0010100101001111,
16'sb0010100110110001,
16'sb0010101000010010,
16'sb0010101001110010,
16'sb0010101011010001,
16'sb0010101100110000,
16'sb0010101110001110,
16'sb0010101111101011,
16'sb0010110001001000,
16'sb0010110010100100,
16'sb0010110100000000,
16'sb0010110101011010,
16'sb0010110110110100,
16'sb0010111000001110,
16'sb0010111001100110,
16'sb0010111010111110,
16'sb0010111100010101,
16'sb0010111101101011,
16'sb0010111111000001,
16'sb0011000000010110,
16'sb0011000001101010,
16'sb0011000010111101,
16'sb0011000100010000,
16'sb0011000101100001,
16'sb0011000110110011,
16'sb0011001000000011,
16'sb0011001001010010,
16'sb0011001010100001,
16'sb0011001011101111,
16'sb0011001100111100,
16'sb0011001110001000,
16'sb0011001111010100,
16'sb0011010000011110,
16'sb0011010001101000,
16'sb0011010010110001,
16'sb0011010011111010,
16'sb0011010101000001,
16'sb0011010110001000,
16'sb0011010111001101,
16'sb0011011000010010,
16'sb0011011001010110,
16'sb0011011010011001,
16'sb0011011011011100,
16'sb0011011100011101,
16'sb0011011101011110,
16'sb0011011110011110,
16'sb0011011111011101,
16'sb0011100000011011,
16'sb0011100001011000,
16'sb0011100010010100,
16'sb0011100011001111,
16'sb0011100100001010,
16'sb0011100101000011,
16'sb0011100101111100,
16'sb0011100110110100,
16'sb0011100111101011,
16'sb0011101000100001,
16'sb0011101001010110,
16'sb0011101010001010,
16'sb0011101010111101,
16'sb0011101011110000,
16'sb0011101100100001,
16'sb0011101101010010,
16'sb0011101110000001,
16'sb0011101110110000,
16'sb0011101111011110,
16'sb0011110000001010,
16'sb0011110000110110,
16'sb0011110001100001,
16'sb0011110010001011,
16'sb0011110010110100,
16'sb0011110011011100,
16'sb0011110100000011,
16'sb0011110100101001,
16'sb0011110101001111,
16'sb0011110101110011,
16'sb0011110110010110,
16'sb0011110110111001,
16'sb0011110111011010,
16'sb0011110111111010,
16'sb0011111000011010,
16'sb0011111000111000,
16'sb0011111001010110,
16'sb0011111001110010,
16'sb0011111010001110,
16'sb0011111010101000,
16'sb0011111011000010,
16'sb0011111011011010,
16'sb0011111011110010,
16'sb0011111100001001,
16'sb0011111100011110,
16'sb0011111100110011,
16'sb0011111101000111,
16'sb0011111101011001,
16'sb0011111101101011,
16'sb0011111101111100,
16'sb0011111110001011,
16'sb0011111110011010,
16'sb0011111110101000,
16'sb0011111110110101,
16'sb0011111111000000,
16'sb0011111111001011,
16'sb0011111111010101,
16'sb0011111111011101,
16'sb0011111111100101,
16'sb0011111111101100,
16'sb0011111111110010,
16'sb0011111111110110,
16'sb0011111111111010,
16'sb0011111111111101,
16'sb0011111111111111,
16'sb0011111111111111,
16'sb0011111111111111,
16'sb0011111111111110,
16'sb0011111111111100,
16'sb0011111111111000,
16'sb0011111111110100,
16'sb0011111111101111,
16'sb0011111111101001,
16'sb0011111111100001,
16'sb0011111111011001,
16'sb0011111111010000,
16'sb0011111111000110,
16'sb0011111110111010,
16'sb0011111110101110,
16'sb0011111110100001,
16'sb0011111110010011,
16'sb0011111110000100,
16'sb0011111101110011,
16'sb0011111101100010,
16'sb0011111101010000,
16'sb0011111100111101,
16'sb0011111100101001,
16'sb0011111100010011,
16'sb0011111011111101,
16'sb0011111011100110,
16'sb0011111011001110,
16'sb0011111010110101,
16'sb0011111010011011,
16'sb0011111010000000,
16'sb0011111001100100,
16'sb0011111001000111,
16'sb0011111000101001,
16'sb0011111000001010,
16'sb0011110111101010,
16'sb0011110111001001,
16'sb0011110110100111,
16'sb0011110110000101,
16'sb0011110101100001,
16'sb0011110100111100,
16'sb0011110100010110,
16'sb0011110011110000,
16'sb0011110011001000,
16'sb0011110010100000,
16'sb0011110001110110,
16'sb0011110001001100,
16'sb0011110000100000,
16'sb0011101111110100,
16'sb0011101111000111,
16'sb0011101110011001,
16'sb0011101101101001,
16'sb0011101100111001,
16'sb0011101100001000,
16'sb0011101011010110,
16'sb0011101010100100,
16'sb0011101001110000,
16'sb0011101000111011,
16'sb0011101000000110,
16'sb0011100111001111,
16'sb0011100110011000,
16'sb0011100101100000,
16'sb0011100100100111,
16'sb0011100011101100,
16'sb0011100010110010,
16'sb0011100001110110,
16'sb0011100000111001,
16'sb0011011111111011,
16'sb0011011110111101,
16'sb0011011101111110,
16'sb0011011100111101,
16'sb0011011011111100,
16'sb0011011010111010,
16'sb0011011001111000,
16'sb0011011000110100,
16'sb0011010111110000,
16'sb0011010110101010,
16'sb0011010101100100,
16'sb0011010100011101,
16'sb0011010011010101,
16'sb0011010010001101,
16'sb0011010001000011,
16'sb0011001111111001,
16'sb0011001110101110,
16'sb0011001101100010,
16'sb0011001100010101,
16'sb0011001011001000,
16'sb0011001001111001,
16'sb0011001000101010,
16'sb0011000111011010,
16'sb0011000110001010,
16'sb0011000100111000,
16'sb0011000011100110,
16'sb0011000010010011,
16'sb0011000000111111,
16'sb0010111111101011,
16'sb0010111110010110,
16'sb0010111101000000,
16'sb0010111011101001,
16'sb0010111010010010,
16'sb0010111000111001,
16'sb0010110111100001,
16'sb0010110110000111,
16'sb0010110100101101,
16'sb0010110011010010,
16'sb0010110001110110,
16'sb0010110000011010,
16'sb0010101110111100,
16'sb0010101101011111,
16'sb0010101100000000,
16'sb0010101010100001,
16'sb0010101001000001,
16'sb0010100111100001,
16'sb0010100110000000,
16'sb0010100100011110,
16'sb0010100010111100,
16'sb0010100001011000,
16'sb0010011111110101,
16'sb0010011110010000,
16'sb0010011100101100,
16'sb0010011011000110,
16'sb0010011001100000,
16'sb0010010111111001,
16'sb0010010110010010,
16'sb0010010100101010,
16'sb0010010011000001,
16'sb0010010001011000,
16'sb0010001111101111,
16'sb0010001110000101,
16'sb0010001100011010,
16'sb0010001010101110,
16'sb0010001001000011,
16'sb0010000111010110,
16'sb0010000101101001,
16'sb0010000011111100,
16'sb0010000010001110,
16'sb0010000000100000,
16'sb0001111110110001,
16'sb0001111101000001,
16'sb0001111011010001,
16'sb0001111001100001,
16'sb0001110111110000,
16'sb0001110101111110,
16'sb0001110100001101,
16'sb0001110010011010,
16'sb0001110000101000,
16'sb0001101110110100,
16'sb0001101101000001,
16'sb0001101011001101,
16'sb0001101001011000,
16'sb0001100111100100,
16'sb0001100101101110,
16'sb0001100011111001,
16'sb0001100010000011,
16'sb0001100000001100,
16'sb0001011110010101,
16'sb0001011100011110,
16'sb0001011010100111,
16'sb0001011000101111,
16'sb0001010110110111,
16'sb0001010100111110,
16'sb0001010011000101,
16'sb0001010001001100,
16'sb0001001111010010,
16'sb0001001101011000,
16'sb0001001011011110,
16'sb0001001001100100,
16'sb0001000111101001,
16'sb0001000101101110,
16'sb0001000011110011,
16'sb0001000001110111,
16'sb0000111111111011,
16'sb0000111101111111,
16'sb0000111100000011,
16'sb0000111010000110,
16'sb0000111000001010,
16'sb0000110110001101,
16'sb0000110100001111,
16'sb0000110010010010,
16'sb0000110000010100,
16'sb0000101110010111,
16'sb0000101100011001,
16'sb0000101010011011,
16'sb0000101000011100,
16'sb0000100110011110,
16'sb0000100100011111,
16'sb0000100010100000,
16'sb0000100000100001,
16'sb0000011110100010,
16'sb0000011100100011,
16'sb0000011010100100,
16'sb0000011000100101,
16'sb0000010110100101,
16'sb0000010100100110,
16'sb0000010010100110,
16'sb0000010000100110,
16'sb0000001110100111,
16'sb0000001100100111,
16'sb0000001010100111,
16'sb0000001000100111,
16'sb0000000110100111,
16'sb0000000100100111,
16'sb0000000010100111,
16'sb0000000000100111,
16'sb1111111110100111,
16'sb1111111100100111,
16'sb1111111010100111,
16'sb1111111000100111,
16'sb1111110110100111,
16'sb1111110100100111,
16'sb1111110010101000,
16'sb1111110000101000,
16'sb1111101110101000,
16'sb1111101100101000,
16'sb1111101010101001,
16'sb1111101000101001,
16'sb1111100110101010,
16'sb1111100100101010,
16'sb1111100010101011,
16'sb1111100000101100,
16'sb1111011110101101,
16'sb1111011100101110
};

assign out = ROM[theta];

endmodule