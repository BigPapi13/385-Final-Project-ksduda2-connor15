
module cos
(
    input [9:0] theta,     //10 bits of precision, first 3 are integer part
    output [15:0] out
);

parameter [0:9][15:0] ROM = {
16'b1000000000000000,
16'b0111111111111111,
16'b0111111111111100,
16'b0111111111110111,
16'b0111111111110000,
16'b0111111111100111,
16'b0111111111011100,
16'b0111111111001111,
16'b0111111111000000,
16'b0111111110101111,
16'b0111111110011100,
16'b0111111110000111,
16'b0111111101110000,
16'b0111111101010111,
16'b0111111100111100,
16'b0111111100011111,
16'b0111111100000000,
16'b0111111011011111,
16'b0111111010111100,
16'b0111111010010111,
16'b0111111001110000,
16'b0111111001000111,
16'b0111111000011101,
16'b0111110111110000,
16'b0111110111000001,
16'b0111110110010000,
16'b0111110101011110,
16'b0111110100101001,
16'b0111110011110011,
16'b0111110010111010,
16'b0111110010000000,
16'b0111110001000011,
16'b0111110000000101,
16'b0111101111000101,
16'b0111101110000010,
16'b0111101100111110,
16'b0111101011111000,
16'b0111101010110000,
16'b0111101001100110,
16'b0111101000011010,
16'b0111100111001100,
16'b0111100101111101,
16'b0111100100101011,
16'b0111100011011000,
16'b0111100010000010,
16'b0111100000101011,
16'b0111011111010010,
16'b0111011101110111,
16'b0111011100011010,
16'b0111011010111100,
16'b0111011001011011,
16'b0111010111111001,
16'b0111010110010100,
16'b0111010100101110,
16'b0111010011000110,
16'b0111010001011101,
16'b0111001111110001,
16'b0111001110000100,
16'b0111001100010101,
16'b0111001010100100,
16'b0111001000110001,
16'b0111000110111100,
16'b0111000101000110,
16'b0111000011001110,
16'b0111000001010100,
16'b0110111111011001,
16'b0110111101011011,
16'b0110111011011100,
16'b0110111001011011,
16'b0110110111011001,
16'b0110110101010100,
16'b0110110011001110,
16'b0110110001000111,
16'b0110101110111101,
16'b0110101100110010,
16'b0110101010100110,
16'b0110101000010111,
16'b0110100110000111,
16'b0110100011110101,
16'b0110100001100010,
16'b0110011111001101,
16'b0110011100110111,
16'b0110011010011110,
16'b0110011000000101,
16'b0110010101101001,
16'b0110010011001100,
16'b0110010000101110,
16'b0110001110001101,
16'b0110001011101100,
16'b0110001001001001,
16'b0110000110100100,
16'b0110000011111101,
16'b0110000001010110,
16'b0101111110101100,
16'b0101111100000010,
16'b0101111001010101,
16'b0101110110100111,
16'b0101110011111000,
16'b0101110001001000,
16'b0101101110010101,
16'b0101101011100010,
16'b0101101000101101,
16'b0101100101110111,
16'b0101100010111111,
16'b0101100000000110,
16'b0101011101001011,
16'b0101011010001111,
16'b0101010111010010,
16'b0101010100010011,
16'b0101010001010011,
16'b0101001110010010,
16'b0101001011010000,
16'b0101001000001100,
16'b0101000101000111,
16'b0101000010000000,
16'b0100111110111000,
16'b0100111011110000,
16'b0100111000100101,
16'b0100110101011010,
16'b0100110010001110,
16'b0100101111000000,
16'b0100101011110001,
16'b0100101000100001,
16'b0100100101001111,
16'b0100100001111101,
16'b0100011110101001,
16'b0100011011010101,
16'b0100010111111111,
16'b0100010100101000,
16'b0100010001010000,
16'b0100001101110111,
16'b0100001010011101,
16'b0100000111000010,
16'b0100000011100110,
16'b0100000000001001,
16'b0011111100101010,
16'b0011111001001011,
16'b0011110101101011,
16'b0011110010001010,
16'b0011101110101000,
16'b0011101011000101,
16'b0011100111100001,
16'b0011100011111101,
16'b0011100000010111,
16'b0011011100110000,
16'b0011011001001001,
16'b0011010101100001,
16'b0011010001111000,
16'b0011001110001110,
16'b0011001010100011,
16'b0011000110110111,
16'b0011000011001011,
16'b0010111111011110,
16'b0010111011110000,
16'b0010111000000010,
16'b0010110100010010,
16'b0010110000100011,
16'b0010101100110010,
16'b0010101001000001,
16'b0010100101001111,
16'b0010100001011100,
16'b0010011101101001,
16'b0010011001110101,
16'b0010010110000000,
16'b0010010010001011,
16'b0010001110010110,
16'b0010001010100000,
16'b0010000110101001,
16'b0010000010110010,
16'b0001111110111010,
16'b0001111011000010,
16'b0001110111001001,
16'b0001110011010000,
16'b0001101111010110,
16'b0001101011011100,
16'b0001100111100001,
16'b0001100011100110,
16'b0001011111101011,
16'b0001011011101111,
16'b0001010111110011,
16'b0001010011110111,
16'b0001001111111010,
16'b0001001011111101,
16'b0001001000000000,
16'b0001000100000010,
16'b0001000000000101,
16'b0000111100000110,
16'b0000111000001000,
16'b0000110100001010,
16'b0000110000001011,
16'b0000101100001100,
16'b0000101000001101,
16'b0000100100001101,
16'b0000100000001110,
16'b0000011100001110,
16'b0000011000001111,
16'b0000010100001111,
16'b0000010000001111,
16'b0000001100001111,
16'b0000001000001111,
16'b0000000100001111,
16'b0000000000001111,
16'b1111111100001111,
16'b1111111000001111,
16'b1111110100001111,
16'b1111110000010000,
16'b1111101100010000,
16'b1111101000010000,
16'b1111100100010000,
16'b1111100000010001,
16'b1111011100010001,
16'b1111011000010010,
16'b1111010100010011,
16'b1111010000010100,
16'b1111001100010101,
16'b1111001000010110,
16'b1111000100011000,
16'b1111000000011010,
16'b1110111100011100,
16'b1110111000011110,
16'b1110110100100001,
16'b1110110000100100,
16'b1110101100100111,
16'b1110101000101011,
16'b1110100100101111,
16'b1110100000110011,
16'b1110011100111000,
16'b1110011000111101,
16'b1110010101000010,
16'b1110010001001000,
16'b1110001101001110,
16'b1110001001010101,
16'b1110000101011100,
16'b1110000001100100,
16'b1101111101101100,
16'b1101111001110101,
16'b1101110101111110,
16'b1101110010001000,
16'b1101101110010010,
16'b1101101010011101,
16'b1101100110101000,
16'b1101100010110100,
16'b1101011111000001,
16'b1101011011001110,
16'b1101010111011100,
16'b1101010011101011,
16'b1101001111111010,
16'b1101001100001010,
16'b1101001000011011,
16'b1101000100101100,
16'b1101000000111110,
16'b1100111101010001,
16'b1100111001100101,
16'b1100110101111001,
16'b1100110010001110,
16'b1100101110100100,
16'b1100101010111011,
16'b1100100111010011,
16'b1100100011101011,
16'b1100100000000101,
16'b1100011100011111,
16'b1100011000111010,
16'b1100010101010110,
16'b1100010001110011,
16'b1100001110010001,
16'b1100001010110000,
16'b1100000111001111,
16'b1100000011110000,
16'b1100000000010010,
16'b1011111100110101,
16'b1011111001011000,
16'b1011110101111101,
16'b1011110010100011,
16'b1011101111001010,
16'b1011101011110010,
16'b1011101000011011,
16'b1011100101000101,
16'b1011100001110000,
16'b1011011110011100,
16'b1011011011001010,
16'b1011010111111000,
16'b1011010100101000,
16'b1011010001011001,
16'b1011001110001011,
16'b1011001010111110,
16'b1011000111110011,
16'b1011000100101000,
16'b1011000001011111,
16'b1010111110011000,
16'b1010111011010001,
16'b1010111000001100,
16'b1010110101001000,
16'b1010110010000101,
16'b1010101111000100,
16'b1010101100000011,
16'b1010101001000101,
16'b1010100110000111,
16'b1010100011001011,
16'b1010100000010000,
16'b1010011101010111,
16'b1010011010011111,
16'b1010010111101001,
16'b1010010100110011,
16'b1010010010000000,
16'b1010001111001101,
16'b1010001100011101,
16'b1010001001101101,
16'b1010000110111111,
16'b1010000100010011,
16'b1010000001101000,
16'b1001111110111110,
16'b1001111100010110,
16'b1001111001110000,
16'b1001110111001011,
16'b1001110100100111,
16'b1001110010000110,
16'b1001101111100101,
16'b1001101101000110,
16'b1001101010101001,
16'b1001101000001110,
16'b1001100101110100,
16'b1001100011011011,
16'b1001100001000100,
16'b1001011110101111,
16'b1001011100011100,
16'b1001011010001010,
16'b1001010111111010,
16'b1001010101101011,
16'b1001010011011110,
16'b1001010001010011,
16'b1001001111001001,
16'b1001001101000001,
16'b1001001010111011,
16'b1001001000110111,
16'b1001000110110100,
16'b1001000100110011,
16'b1001000010110011,
16'b1001000000110110,
16'b1000111110111010,
16'b1000111101000000,
16'b1000111011001000,
16'b1000111001010001,
16'b1000110111011100,
16'b1000110101101001,
16'b1000110011111000,
16'b1000110010001001,
16'b1000110000011011,
16'b1000101110101111,
16'b1000101101000110,
16'b1000101011011101,
16'b1000101001110111,
16'b1000101000010011,
16'b1000100110110000,
16'b1000100101001111,
16'b1000100011110000,
16'b1000100010010011,
16'b1000100000111000,
16'b1000011111011111,
16'b1000011110000111,
16'b1000011100110010,
16'b1000011011011110,
16'b1000011010001100,
16'b1000011000111100,
16'b1000010111101110,
16'b1000010110100010,
16'b1000010101011000,
16'b1000010100010000,
16'b1000010011001001,
16'b1000010010000101,
16'b1000010001000011,
16'b1000010000000010,
16'b1000001111000011,
16'b1000001110000111,
16'b1000001101001100,
16'b1000001100010011,
16'b1000001011011100,
16'b1000001010101000,
16'b1000001001110101,
16'b1000001001000100,
16'b1000001000010101,
16'b1000000111101000,
16'b1000000110111101,
16'b1000000110010100,
16'b1000000101101101,
16'b1000000101000111,
16'b1000000100100100,
16'b1000000100000011,
16'b1000000011100100,
16'b1000000011000111,
16'b1000000010101100,
16'b1000000010010010,
16'b1000000001111011,
16'b1000000001100110,
16'b1000000001010011,
16'b1000000001000001,
16'b1000000000110010,
16'b1000000000100101,
16'b1000000000011010,
16'b1000000000010001,
16'b1000000000001001,
16'b1000000000000100,
16'b1000000000000001,
16'b1000000000000000,
16'b1000000000000000,
16'b1000000000000011,
16'b1000000000001000,
16'b1000000000001111,
16'b1000000000010111,
16'b1000000000100010,
16'b1000000000101111,
16'b1000000000111110,
16'b1000000001001110,
16'b1000000001100001,
16'b1000000001110110,
16'b1000000010001100,
16'b1000000010100101,
16'b1000000011000000,
16'b1000000011011101,
16'b1000000011111011,
16'b1000000100011100,
16'b1000000100111111,
16'b1000000101100011,
16'b1000000110001010,
16'b1000000110110010,
16'b1000000111011101,
16'b1000001000001001,
16'b1000001000111000,
16'b1000001001101000,
16'b1000001010011011,
16'b1000001011001111,
16'b1000001100000110,
16'b1000001100111110,
16'b1000001101111000,
16'b1000001110110100,
16'b1000001111110010,
16'b1000010000110010,
16'b1000010001110100,
16'b1000010010111000,
16'b1000010011111110,
16'b1000010101000110,
16'b1000010110010000,
16'b1000010111011011,
16'b1000011000101001,
16'b1000011001111000,
16'b1000011011001010,
16'b1000011100011101,
16'b1000011101110010,
16'b1000011111001001,
16'b1000100000100010,
16'b1000100001111100,
16'b1000100011011001,
16'b1000100100110111,
16'b1000100110011000,
16'b1000100111111010,
16'b1000101001011110,
16'b1000101011000100,
16'b1000101100101100,
16'b1000101110010101,
16'b1000110000000000,
16'b1000110001101110,
16'b1000110011011100,
16'b1000110101001101,
16'b1000110111000000,
16'b1000111000110100,
16'b1000111010101010,
16'b1000111100100010,
16'b1000111110011100,
16'b1001000000010111,
16'b1001000010010100,
16'b1001000100010011,
16'b1001000110010100,
16'b1001001000010110,
16'b1001001010011010,
16'b1001001100100000,
16'b1001001110100111,
16'b1001010000110001,
16'b1001010010111011,
16'b1001010101001000,
16'b1001010111010110,
16'b1001011001100110,
16'b1001011011110111,
16'b1001011110001011,
16'b1001100000011111,
16'b1001100010110110,
16'b1001100101001110,
16'b1001100111100111,
16'b1001101010000011,
16'b1001101100011111,
16'b1001101110111110,
16'b1001110001011110,
16'b1001110011111111,
16'b1001110110100010,
16'b1001111001000111,
16'b1001111011101101,
16'b1001111110010100,
16'b1010000000111110,
16'b1010000011101000,
16'b1010000110010100,
16'b1010001001000010,
16'b1010001011110001,
16'b1010001110100001,
16'b1010010001010011,
16'b1010010100000111,
16'b1010010110111100,
16'b1010011001110010,
16'b1010011100101001,
16'b1010011111100010,
16'b1010100010011101,
16'b1010100101011001,
16'b1010101000010110,
16'b1010101011010100,
16'b1010101110010100,
16'b1010110001010101,
16'b1010110100010111,
16'b1010110111011011,
16'b1010111010100000,
16'b1010111101100110,
16'b1011000000101110,
16'b1011000011110110,
16'b1011000111000000,
16'b1011001010001100,
16'b1011001101011000,
16'b1011010000100110,
16'b1011010011110100,
16'b1011010111000100,
16'b1011011010010110,
16'b1011011101101000,
16'b1011100000111011,
16'b1011100100010000,
16'b1011100111100101,
16'b1011101010111100,
16'b1011101110010100,
16'b1011110001101101,
16'b1011110101000111,
16'b1011111000100010,
16'b1011111011111110,
16'b1011111111011011,
16'b1100000010111001,
16'b1100000110011000,
16'b1100001001111000,
16'b1100001101011001,
16'b1100010000111011,
16'b1100010100011110,
16'b1100011000000001,
16'b1100011011100110,
16'b1100011111001100,
16'b1100100010110010,
16'b1100100110011001,
16'b1100101010000010,
16'b1100101101101011,
16'b1100110001010100,
16'b1100110100111111,
16'b1100111000101010,
16'b1100111100010111,
16'b1101000000000100,
16'b1101000011110001,
16'b1101000111100000,
16'b1101001011001111,
16'b1101001110111111,
16'b1101010010101111,
16'b1101010110100000,
16'b1101011010010010,
16'b1101011110000101,
16'b1101100001111000,
16'b1101100101101100,
16'b1101101001100000,
16'b1101101101010101,
16'b1101110001001011,
16'b1101110101000001,
16'b1101111000111000,
16'b1101111100101111,
16'b1110000000100110,
16'b1110000100011111,
16'b1110001000010111,
16'b1110001100010001,
16'b1110010000001010,
16'b1110010100000100,
16'b1110010111111111,
16'b1110011011111001,
16'b1110011111110101,
16'b1110100011110000,
16'b1110100111101100,
16'b1110101011101001,
16'b1110101111100101,
16'b1110110011100010,
16'b1110110111100000,
16'b1110111011011101,
16'b1110111111011011,
16'b1111000011011001,
16'b1111000111010111,
16'b1111001011010110,
16'b1111001111010101,
16'b1111010011010100,
16'b1111010111010011,
16'b1111011011010010,
16'b1111011111010001,
16'b1111100011010001,
16'b1111100111010001,
16'b1111101011010000,
16'b1111101111010000,
16'b1111110011010000,
16'b1111110111010000,
16'b1111111011010000,
16'b1111111111010000,
16'b0000000011010000,
16'b0000000111010000,
16'b0000001011010000,
16'b0000001111010000,
16'b0000010011010000,
16'b0000010111001111,
16'b0000011011001111,
16'b0000011111001111,
16'b0000100011001110,
16'b0000100111001101,
16'b0000101011001101,
16'b0000101111001100,
16'b0000110011001010,
16'b0000110111001001,
16'b0000111011000111,
16'b0000111111000110,
16'b0001000011000100,
16'b0001000111000001,
16'b0001001010111111,
16'b0001001110111100,
16'b0001010010111000,
16'b0001010110110101,
16'b0001011010110001,
16'b0001011110101101,
16'b0001100010101000,
16'b0001100110100011,
16'b0001101010011110,
16'b0001101110011000,
16'b0001110010010010,
16'b0001110110001011,
16'b0001111010000100,
16'b0001111101111100,
16'b0010000001110100,
16'b0010000101101100,
16'b0010001001100010,
16'b0010001101011001,
16'b0010010001001111,
16'b0010010101000100,
16'b0010011000111000,
16'b0010011100101100,
16'b0010100000100000,
16'b0010100100010011,
16'b0010101000000101,
16'b0010101011110110,
16'b0010101111100111,
16'b0010110011010111,
16'b0010110111000111,
16'b0010111010110101,
16'b0010111110100011,
16'b0011000010010000,
16'b0011000101111101,
16'b0011001001101001,
16'b0011001101010100,
16'b0011010000111110,
16'b0011010100100111,
16'b0011011000001111,
16'b0011011011110111,
16'b0011011111011110,
16'b0011100011000100,
16'b0011100110101001,
16'b0011101010001101,
16'b0011101101110000,
16'b0011110001010010,
16'b0011110100110100,
16'b0011111000010100,
16'b0011111011110011,
16'b0011111111010010,
16'b0100000010101111,
16'b0100000110001100,
16'b0100001001100111,
16'b0100001101000001,
16'b0100010000011011,
16'b0100010011110011,
16'b0100010111001010,
16'b0100011010100000,
16'b0100011101110101,
16'b0100100001001001,
16'b0100100100011011,
16'b0100100111101101,
16'b0100101010111101,
16'b0100101110001101,
16'b0100110001011011,
16'b0100110100101000,
16'b0100110111110011,
16'b0100111010111110,
16'b0100111110000111,
16'b0101000001001111,
16'b0101000100010110,
16'b0101000111011011,
16'b0101001010011111,
16'b0101001101100010,
16'b0101010000100100,
16'b0101010011100100,
16'b0101010110100011,
16'b0101011001100000,
16'b0101011100011101,
16'b0101011111010111,
16'b0101100010010001,
16'b0101100101001001,
16'b0101101000000000,
16'b0101101010110101,
16'b0101101101101001,
16'b0101110000011100,
16'b0101110011001101,
16'b0101110101111100,
16'b0101111000101010,
16'b0101111011010111,
16'b0101111110000010,
16'b0110000000101100,
16'b0110000011010100,
16'b0110000101111011,
16'b0110001000100000,
16'b0110001011000011,
16'b0110001101100110,
16'b0110010000000110,
16'b0110010010100101,
16'b0110010101000010,
16'b0110010111011110,
16'b0110011001111000,
16'b0110011100010001,
16'b0110011110101000,
16'b0110100000111101,
16'b0110100011010001,
16'b0110100101100011,
16'b0110100111110100,
16'b0110101010000010,
16'b0110101100010000,
16'b0110101110011011,
16'b0110110000100101,
16'b0110110010101101,
16'b0110110100110011,
16'b0110110110111000,
16'b0110111000111011,
16'b0110111010111100,
16'b0110111100111100,
16'b0110111110111010,
16'b0111000000110110,
16'b0111000010110000,
16'b0111000100101000,
16'b0111000110011111,
16'b0111001000010100,
16'b0111001010000111,
16'b0111001011111001,
16'b0111001101101000,
16'b0111001111010110,
16'b0111010001000010,
16'b0111010010101100,
16'b0111010100010101,
16'b0111010101111011,
16'b0111010111100000,
16'b0111011001000011,
16'b0111011010100100,
16'b0111011100000011,
16'b0111011101100000,
16'b0111011110111100,
16'b0111100000010101,
16'b0111100001101101,
16'b0111100011000011,
16'b0111100100010111,
16'b0111100101101001,
16'b0111100110111001,
16'b0111101000000111,
16'b0111101001010011,
16'b0111101010011110,
16'b0111101011100110,
16'b0111101100101101,
16'b0111101101110010,
16'b0111101110110100,
16'b0111101111110101,
16'b0111110000110100,
16'b0111110001110001,
16'b0111110010101100,
16'b0111110011100101,
16'b0111110100011100,
16'b0111110101010001,
16'b0111110110000100,
16'b0111110110110101,
16'b0111110111100101,
16'b0111111000010010,
16'b0111111000111101,
16'b0111111001100110,
16'b0111111010001110,
16'b0111111010110011,
16'b0111111011010110,
16'b0111111011111000,
16'b0111111100010111,
16'b0111111100110101,
16'b0111111101010000,
16'b0111111101101010,
16'b0111111110000001,
16'b0111111110010111,
16'b0111111110101010,
16'b0111111110111011,
16'b0111111111001011,
16'b0111111111011000,
16'b0111111111100100,
16'b0111111111101101,
16'b0111111111110101,
16'b0111111111111010,
16'b0111111111111110,
16'b0111111111111111,
16'b0111111111111111,
16'b0111111111111100,
16'b0111111111111000,
16'b0111111111110001,
16'b0111111111101001,
16'b0111111111011110,
16'b0111111111010010,
16'b0111111111000011,
16'b0111111110110011,
16'b0111111110100000,
16'b0111111110001100,
16'b0111111101110101,
16'b0111111101011101,
16'b0111111101000011,
16'b0111111100100110,
16'b0111111100001000,
16'b0111111011100111,
16'b0111111011000101,
16'b0111111010100000,
16'b0111111001111010,
16'b0111111001010010,
16'b0111111000100111,
16'b0111110111111011,
16'b0111110111001101,
16'b0111110110011101,
16'b0111110101101011,
16'b0111110100110110,
16'b0111110100000000,
16'b0111110011001000,
16'b0111110010001110,
16'b0111110001010010,
16'b0111110000010100,
16'b0111101111010101,
16'b0111101110010011,
16'b0111101101001111,
16'b0111101100001010,
16'b0111101011000010,
16'b0111101001111001,
16'b0111101000101101,
16'b0111100111100000,
16'b0111100110010001,
16'b0111100101000000,
16'b0111100011101101,
16'b0111100010011000,
16'b0111100001000001,
16'b0111011111101000,
16'b0111011110001110,
16'b0111011100110010,
16'b0111011011010011,
16'b0111011001110011,
16'b0111011000010001,
16'b0111010110101101,
16'b0111010101001000,
16'b0111010011100000,
16'b0111010001110111,
16'b0111010000001100,
16'b0111001110011111,
16'b0111001100110000,
16'b0111001011000000,
16'b0111001001001110,
16'b0111000111011001,
16'b0111000101100100,
16'b0111000011101100,
16'b0111000001110010,
16'b0110111111110111,
16'b0110111101111010,
16'b0110111011111100,
16'b0110111001111011,
16'b0110110111111001,
16'b0110110101110101,
16'b0110110011110000,
16'b0110110001101001,
16'b0110101111100000,
16'b0110101101010101,
16'b0110101011001001,
16'b0110101000111011,
16'b0110100110101011,
16'b0110100100011010,
16'b0110100010000111,
16'b0110011111110010,
16'b0110011101011100,
16'b0110011011000100,
16'b0110011000101011,
16'b0110010110010000,
16'b0110010011110011,
16'b0110010001010101,
16'b0110001110110101,
16'b0110001100010100,
16'b0110001001110001,
16'b0110000111001101,
16'b0110000100100111,
16'b0110000001111111,
16'b0101111111010110,
16'b0101111100101100,
16'b0101111010000000,
16'b0101110111010011,
16'b0101110100100100,
16'b0101110001110011,
16'b0101101111000010,
16'b0101101100001111,
16'b0101101001011010,
16'b0101100110100100,
16'b0101100011101100,
16'b0101100000110100,
16'b0101011101111001,
16'b0101011010111110,
16'b0101011000000001,
16'b0101010101000011,
16'b0101010010000011,
16'b0101001111000010,
16'b0101001100000000,
16'b0101001000111100,
16'b0101000101111000,
16'b0101000010110001,
16'b0100111111101010,
16'b0100111100100001,
16'b0100111001011000,
16'b0100110110001101,
16'b0100110011000000,
16'b0100101111110011,
16'b0100101100100100,
16'b0100101001010100,
16'b0100100110000011,
16'b0100100010110001,
16'b0100011111011110,
16'b0100011100001010,
16'b0100011000110100,
16'b0100010101011101,
16'b0100010010000110,
16'b0100001110101101,
16'b0100001011010011,
16'b0100000111111000,
16'b0100000100011100,
16'b0100000001000000,
16'b0011111101100010,
16'b0011111010000011,
16'b0011110110100011,
16'b0011110011000010,
16'b0011101111100000,
16'b0011101011111101,
16'b0011101000011010,
16'b0011100100110101,
16'b0011100001010000,
16'b0011011101101001,
16'b0011011010000010,
16'b0011010110011010,
16'b0011010010110001,
16'b0011001111001000,
16'b0011001011011101,
16'b0011000111110010,
16'b0011000100000110,
16'b0011000000011001,
16'b0010111100101011,
16'b0010111000111101,
16'b0010110101001110,
16'b0010110001011110,
16'b0010101101101110,
16'b0010101001111100,
16'b0010100110001011,
16'b0010100010011000,
16'b0010011110100101,
16'b0010011010110001,
16'b0010010110111101,
16'b0010010011001000,
16'b0010001111010011,
16'b0010001011011101,
16'b0010000111100110,
16'b0010000011101111,
16'b0001111111110111,
16'b0001111011111111,
16'b0001111000000110,
16'b0001110100001101,
16'b0001110000010100,
16'b0001101100011010,
16'b0001101000011111,
16'b0001100100100101,
16'b0001100000101001,
16'b0001011100101110,
16'b0001011000110010,
16'b0001010100110110,
16'b0001010000111001,
16'b0001001100111100,
16'b0001001000111111,
16'b0001000101000001,
16'b0001000001000011,
16'b0000111101000101,
16'b0000111001000111,
16'b0000110101001001,
16'b0000110001001010,
16'b0000101101001011,
16'b0000101001001100,
16'b0000100101001101,
16'b0000100001001101,
16'b0000011101001110,
16'b0000011001001110,
16'b0000010101001110,
16'b0000010001001111,
16'b0000001101001111,
16'b0000001001001111,
16'b0000000101001111,
16'b0000000001001111,
16'b1111111101001111,
16'b1111111001001111,
16'b1111110101001111,
16'b1111110001001111,
16'b1111101101001111,
16'b1111101001001111,
16'b1111100101010000,
16'b1111100001010000,
16'b1111011101010000,
16'b1111011001010001,
16'b1111010101010010,
16'b1111010001010011,
16'b1111001101010100,
16'b1111001001010101,
16'b1111000101010111,
16'b1111000001011001,
16'b1110111101011011,
16'b1110111001011101
};

assign out = ROM[theta];

endmodule