
// Parameters

module obb_reg
(
    output logic signed [7 : 0] width,
    output logic signed [7 : 0] height,
    output logic signed [31 : 0] pos [1 : 0],
    output logic signed [31 : 0] vel [1 : 0],
    output logic signed [9 : 0] angle
);

always_comb begin


end

endmodule