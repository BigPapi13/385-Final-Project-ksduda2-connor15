
module sin
(
    input [9:0] theta,     //10 bits of precision, first 3 are integer part
    output [15:0] out
);

parameter [0:9][15:0] ROM = {
16'b0000000000000000,
16'b0000000011111111,
16'b0000000111111111,
16'b0000001011111111,
16'b0000001111111111,
16'b0000010011111111,
16'b0000010111111111,
16'b0000011011111111,
16'b0000011111111110,
16'b0000100011111110,
16'b0000100111111101,
16'b0000101011111100,
16'b0000101111111011,
16'b0000110011111010,
16'b0000110111111000,
16'b0000111011110111,
16'b0000111111110101,
16'b0001000011110011,
16'b0001000111110000,
16'b0001001011101110,
16'b0001001111101011,
16'b0001010011100111,
16'b0001010111100100,
16'b0001011011100000,
16'b0001011111011100,
16'b0001100011010111,
16'b0001100111010010,
16'b0001101011001100,
16'b0001101111000110,
16'b0001110011000000,
16'b0001110110111001,
16'b0001111010110010,
16'b0001111110101010,
16'b0010000010100010,
16'b0010000110011010,
16'b0010001010010000,
16'b0010001110000110,
16'b0010010001111100,
16'b0010010101110001,
16'b0010011001100110,
16'b0010011101011010,
16'b0010100001001101,
16'b0010100101000000,
16'b0010101000110010,
16'b0010101100100011,
16'b0010110000010100,
16'b0010110100000100,
16'b0010110111110011,
16'b0010111011100010,
16'b0010111111001111,
16'b0011000010111100,
16'b0011000110101001,
16'b0011001010010100,
16'b0011001101111111,
16'b0011010001101001,
16'b0011010101010010,
16'b0011011000111011,
16'b0011011100100010,
16'b0011100000001001,
16'b0011100011101110,
16'b0011100111010011,
16'b0011101010110111,
16'b0011101110011010,
16'b0011110001111100,
16'b0011110101011101,
16'b0011111000111101,
16'b0011111100011101,
16'b0011111111111011,
16'b0100000011011000,
16'b0100000110110100,
16'b0100001010010000,
16'b0100001101101010,
16'b0100010001000011,
16'b0100010100011011,
16'b0100010111110010,
16'b0100011011001000,
16'b0100011110011100,
16'b0100100001110000,
16'b0100100101000010,
16'b0100101000010100,
16'b0100101011100100,
16'b0100101110110011,
16'b0100110010000001,
16'b0100110101001101,
16'b0100111000011001,
16'b0100111011100011,
16'b0100111110101100,
16'b0101000001110100,
16'b0101000100111010,
16'b0101001000000000,
16'b0101001011000011,
16'b0101001110000110,
16'b0101010001000111,
16'b0101010100000111,
16'b0101010111000110,
16'b0101011010000011,
16'b0101011100111111,
16'b0101011111111010,
16'b0101100010110011,
16'b0101100101101011,
16'b0101101000100010,
16'b0101101011010111,
16'b0101101110001010,
16'b0101110000111101,
16'b0101110011101101,
16'b0101110110011101,
16'b0101111001001011,
16'b0101111011110111,
16'b0101111110100010,
16'b0110000001001011,
16'b0110000011110011,
16'b0110000110011010,
16'b0110001000111110,
16'b0110001011100010,
16'b0110001110000011,
16'b0110010000100100,
16'b0110010011000010,
16'b0110010101011111,
16'b0110010111111011,
16'b0110011010010101,
16'b0110011100101101,
16'b0110011111000100,
16'b0110100001011001,
16'b0110100011101100,
16'b0110100101111110,
16'b0110101000001110,
16'b0110101010011101,
16'b0110101100101010,
16'b0110101110110101,
16'b0110110000111110,
16'b0110110011000110,
16'b0110110101001100,
16'b0110110111010001,
16'b0110111001010011,
16'b0110111011010100,
16'b0110111101010011,
16'b0110111111010001,
16'b0111000001001101,
16'b0111000011000110,
16'b0111000100111111,
16'b0111000110110101,
16'b0111001000101010,
16'b0111001010011101,
16'b0111001100001110,
16'b0111001101111101,
16'b0111001111101010,
16'b0111010001010110,
16'b0111010011000000,
16'b0111010100101000,
16'b0111010110001110,
16'b0111010111110011,
16'b0111011001010101,
16'b0111011010110110,
16'b0111011100010101,
16'b0111011101110010,
16'b0111011111001101,
16'b0111100000100110,
16'b0111100001111101,
16'b0111100011010011,
16'b0111100100100110,
16'b0111100101111000,
16'b0111100111001000,
16'b0111101000010101,
16'b0111101001100001,
16'b0111101010101011,
16'b0111101011110100,
16'b0111101100111010,
16'b0111101101111110,
16'b0111101111000000,
16'b0111110000000001,
16'b0111110000111111,
16'b0111110001111100,
16'b0111110010110111,
16'b0111110011101111,
16'b0111110100100110,
16'b0111110101011011,
16'b0111110110001101,
16'b0111110110111110,
16'b0111110111101101,
16'b0111111000011010,
16'b0111111001000101,
16'b0111111001101110,
16'b0111111010010101,
16'b0111111010111010,
16'b0111111011011101,
16'b0111111011111110,
16'b0111111100011101,
16'b0111111100111010,
16'b0111111101010101,
16'b0111111101101110,
16'b0111111110000101,
16'b0111111110011010,
16'b0111111110101101,
16'b0111111110111111,
16'b0111111111001110,
16'b0111111111011011,
16'b0111111111100110,
16'b0111111111101111,
16'b0111111111110110,
16'b0111111111111011,
16'b0111111111111110,
16'b0111111111111111,
16'b0111111111111111,
16'b0111111111111100,
16'b0111111111110111,
16'b0111111111110000,
16'b0111111111100111,
16'b0111111111011100,
16'b0111111111001111,
16'b0111111111000001,
16'b0111111110110000,
16'b0111111110011101,
16'b0111111110001000,
16'b0111111101110001,
16'b0111111101011000,
16'b0111111100111101,
16'b0111111100100001,
16'b0111111100000010,
16'b0111111011100001,
16'b0111111010111110,
16'b0111111010011010,
16'b0111111001110011,
16'b0111111001001010,
16'b0111111000011111,
16'b0111110111110011,
16'b0111110111000100,
16'b0111110110010100,
16'b0111110101100001,
16'b0111110100101101,
16'b0111110011110110,
16'b0111110010111110,
16'b0111110010000011,
16'b0111110001000111,
16'b0111110000001001,
16'b0111101111001001,
16'b0111101110000110,
16'b0111101101000010,
16'b0111101011111100,
16'b0111101010110101,
16'b0111101001101011,
16'b0111101000011111,
16'b0111100111010001,
16'b0111100110000010,
16'b0111100100110000,
16'b0111100011011101,
16'b0111100010001000,
16'b0111100000110001,
16'b0111011111011000,
16'b0111011101111101,
16'b0111011100100000,
16'b0111011011000010,
16'b0111011001100001,
16'b0111010111111111,
16'b0111010110011011,
16'b0111010100110101,
16'b0111010011001101,
16'b0111010001100011,
16'b0111001111111000,
16'b0111001110001011,
16'b0111001100011100,
16'b0111001010101011,
16'b0111001000111000,
16'b0111000111000100,
16'b0111000101001101,
16'b0111000011010101,
16'b0111000001011100,
16'b0110111111100000,
16'b0110111101100011,
16'b0110111011100100,
16'b0110111001100011,
16'b0110110111100001,
16'b0110110101011101,
16'b0110110011010111,
16'b0110110001001111,
16'b0110101111000110,
16'b0110101100111011,
16'b0110101010101110,
16'b0110101000100000,
16'b0110100110010000,
16'b0110100011111111,
16'b0110100001101011,
16'b0110011111010110,
16'b0110011101000000,
16'b0110011010101000,
16'b0110011000001110,
16'b0110010101110011,
16'b0110010011010110,
16'b0110010000110111,
16'b0110001110010111,
16'b0110001011110110,
16'b0110001001010011,
16'b0110000110101110,
16'b0110000100001000,
16'b0110000001100000,
16'b0101111110110111,
16'b0101111100001100,
16'b0101111001100000,
16'b0101110110110010,
16'b0101110100000011,
16'b0101110001010011,
16'b0101101110100001,
16'b0101101011101101,
16'b0101101000111000,
16'b0101100110000010,
16'b0101100011001010,
16'b0101100000010001,
16'b0101011101010111,
16'b0101011010011011,
16'b0101010111011110,
16'b0101010100011111,
16'b0101010001011111,
16'b0101001110011110,
16'b0101001011011100,
16'b0101001000011000,
16'b0101000101010011,
16'b0101000010001100,
16'b0100111111000101,
16'b0100111011111100,
16'b0100111000110010,
16'b0100110101100111,
16'b0100110010011010,
16'b0100101111001101,
16'b0100101011111110,
16'b0100101000101110,
16'b0100100101011100,
16'b0100100010001010,
16'b0100011110110111,
16'b0100011011100010,
16'b0100011000001100,
16'b0100010100110101,
16'b0100010001011110,
16'b0100001110000101,
16'b0100001010101011,
16'b0100000111010000,
16'b0100000011110011,
16'b0100000000010110,
16'b0011111100111000,
16'b0011111001011001,
16'b0011110101111001,
16'b0011110010011000,
16'b0011101110110110,
16'b0011101011010011,
16'b0011100111101111,
16'b0011100100001011,
16'b0011100000100101,
16'b0011011100111111,
16'b0011011001010111,
16'b0011010101101111,
16'b0011010010000110,
16'b0011001110011100,
16'b0011001010110001,
16'b0011000111000110,
16'b0011000011011010,
16'b0010111111101101,
16'b0010111011111111,
16'b0010111000010001,
16'b0010110100100001,
16'b0010110000110001,
16'b0010101101000001,
16'b0010101001010000,
16'b0010100101011110,
16'b0010100001101011,
16'b0010011101111000,
16'b0010011010000100,
16'b0010010110010000,
16'b0010010010011011,
16'b0010001110100101,
16'b0010001010101111,
16'b0010000110111000,
16'b0010000011000001,
16'b0001111111001001,
16'b0001111011010001,
16'b0001110111011000,
16'b0001110011011111,
16'b0001101111100101,
16'b0001101011101011,
16'b0001100111110001,
16'b0001100011110110,
16'b0001011111111011,
16'b0001011011111111,
16'b0001011000000011,
16'b0001010100000111,
16'b0001010000001010,
16'b0001001100001101,
16'b0001001000010000,
16'b0001000100010010,
16'b0001000000010100,
16'b0000111100010110,
16'b0000111000011000,
16'b0000110100011001,
16'b0000110000011011,
16'b0000101100011100,
16'b0000101000011101,
16'b0000100100011101,
16'b0000100000011110,
16'b0000011100011110,
16'b0000011000011111,
16'b0000010100011111,
16'b0000010000011111,
16'b0000001100011111,
16'b0000001000011111,
16'b0000000100011111,
16'b0000000000011111,
16'b1111111100011111,
16'b1111111000011111,
16'b1111110100011111,
16'b1111110000011111,
16'b1111101100100000,
16'b1111101000100000,
16'b1111100100100000,
16'b1111100000100000,
16'b1111011100100001,
16'b1111011000100010,
16'b1111010100100011,
16'b1111010000100100,
16'b1111001100100101,
16'b1111001000100110,
16'b1111000100101000,
16'b1111000000101010,
16'b1110111100101100,
16'b1110111000101110,
16'b1110110100110001,
16'b1110110000110100,
16'b1110101100110111,
16'b1110101000111010,
16'b1110100100111110,
16'b1110100001000011,
16'b1110011101000111,
16'b1110011001001100,
16'b1110010101010010,
16'b1110010001010111,
16'b1110001101011110,
16'b1110001001100100,
16'b1110000101101100,
16'b1110000001110011,
16'b1101111101111011,
16'b1101111010000100,
16'b1101110110001101,
16'b1101110010010111,
16'b1101101110100001,
16'b1101101010101100,
16'b1101100110111000,
16'b1101100011000100,
16'b1101011111010000,
16'b1101011011011101,
16'b1101010111101011,
16'b1101010011111010,
16'b1101010000001001,
16'b1101001100011001,
16'b1101001000101010,
16'b1101000100111011,
16'b1101000001001101,
16'b1100111101100000,
16'b1100111001110011,
16'b1100110110001000,
16'b1100110010011101,
16'b1100101110110011,
16'b1100101011001010,
16'b1100100111100001,
16'b1100100011111010,
16'b1100100000010011,
16'b1100011100101101,
16'b1100011001001000,
16'b1100010101100100,
16'b1100010010000001,
16'b1100001110011111,
16'b1100001010111110,
16'b1100000111011101,
16'b1100000011111110,
16'b1100000000100000,
16'b1011111101000010,
16'b1011111001100110,
16'b1011110110001011,
16'b1011110010110000,
16'b1011101111010111,
16'b1011101011111111,
16'b1011101000101000,
16'b1011100101010010,
16'b1011100001111101,
16'b1011011110101001,
16'b1011011011010111,
16'b1011011000000101,
16'b1011010100110101,
16'b1011010001100110,
16'b1011001110011000,
16'b1011001011001011,
16'b1011000111111111,
16'b1011000100110101,
16'b1011000001101100,
16'b1010111110100100,
16'b1010111011011101,
16'b1010111000011000,
16'b1010110101010100,
16'b1010110010010001,
16'b1010101111001111,
16'b1010101100001111,
16'b1010101001010000,
16'b1010100110010011,
16'b1010100011010111,
16'b1010100000011100,
16'b1010011101100011,
16'b1010011010101011,
16'b1010010111110100,
16'b1010010100111111,
16'b1010010010001011,
16'b1010001111011000,
16'b1010001100100111,
16'b1010001001111000,
16'b1010000111001010,
16'b1010000100011101,
16'b1010000001110010,
16'b1001111111001001,
16'b1001111100100001,
16'b1001111001111010,
16'b1001110111010101,
16'b1001110100110001,
16'b1001110010001111,
16'b1001101111101111,
16'b1001101101010000,
16'b1001101010110011,
16'b1001101000010111,
16'b1001100101111101,
16'b1001100011100101,
16'b1001100001001110,
16'b1001011110111000,
16'b1001011100100101,
16'b1001011010010011,
16'b1001011000000010,
16'b1001010101110100,
16'b1001010011100111,
16'b1001010001011011,
16'b1001001111010010,
16'b1001001101001010,
16'b1001001011000011,
16'b1001001000111111,
16'b1001000110111100,
16'b1001000100111011,
16'b1001000010111011,
16'b1001000000111110,
16'b1000111111000010,
16'b1000111101001000,
16'b1000111011001111,
16'b1000111001011000,
16'b1000110111100100,
16'b1000110101110000,
16'b1000110011111111,
16'b1000110010010000,
16'b1000110000100010,
16'b1000101110110110,
16'b1000101101001100,
16'b1000101011100100,
16'b1000101001111101,
16'b1000101000011001,
16'b1000100110110110,
16'b1000100101010101,
16'b1000100011110110,
16'b1000100010011001,
16'b1000100000111110,
16'b1000011111100100,
16'b1000011110001101,
16'b1000011100110111,
16'b1000011011100011,
16'b1000011010010001,
16'b1000011001000001,
16'b1000010111110011,
16'b1000010110100111,
16'b1000010101011101,
16'b1000010100010100,
16'b1000010011001110,
16'b1000010010001001,
16'b1000010001000111,
16'b1000010000000110,
16'b1000001111000111,
16'b1000001110001010,
16'b1000001101010000,
16'b1000001100010111,
16'b1000001011100000,
16'b1000001010101011,
16'b1000001001111000,
16'b1000001001000111,
16'b1000001000011000,
16'b1000000111101010,
16'b1000000110111111,
16'b1000000110010110,
16'b1000000101101111,
16'b1000000101001010,
16'b1000000100100110,
16'b1000000100000101,
16'b1000000011100110,
16'b1000000011001001,
16'b1000000010101101,
16'b1000000010010100,
16'b1000000001111101,
16'b1000000001100111,
16'b1000000001010100,
16'b1000000001000010,
16'b1000000000110011,
16'b1000000000100110,
16'b1000000000011010,
16'b1000000000010001,
16'b1000000000001010,
16'b1000000000000100,
16'b1000000000000001,
16'b1000000000000000,
16'b1000000000000000,
16'b1000000000000011,
16'b1000000000000111,
16'b1000000000001110,
16'b1000000000010111,
16'b1000000000100001,
16'b1000000000101110,
16'b1000000000111101,
16'b1000000001001101,
16'b1000000001100000,
16'b1000000001110100,
16'b1000000010001011,
16'b1000000010100100,
16'b1000000010111110,
16'b1000000011011011,
16'b1000000011111001,
16'b1000000100011010,
16'b1000000100111100,
16'b1000000101100001,
16'b1000000110000111,
16'b1000000110110000,
16'b1000000111011010,
16'b1000001000000111,
16'b1000001000110101,
16'b1000001001100101,
16'b1000001010011000,
16'b1000001011001100,
16'b1000001100000010,
16'b1000001100111010,
16'b1000001101110100,
16'b1000001110110000,
16'b1000001111101110,
16'b1000010000101110,
16'b1000010001110000,
16'b1000010010110100,
16'b1000010011111010,
16'b1000010101000001,
16'b1000010110001011,
16'b1000010111010111,
16'b1000011000100100,
16'b1000011001110011,
16'b1000011011000100,
16'b1000011100011000,
16'b1000011101101101,
16'b1000011111000011,
16'b1000100000011100,
16'b1000100001110111,
16'b1000100011010011,
16'b1000100100110010,
16'b1000100110010010,
16'b1000100111110100,
16'b1000101001011000,
16'b1000101010111101,
16'b1000101100100101,
16'b1000101110001110,
16'b1000101111111010,
16'b1000110001100111,
16'b1000110011010110,
16'b1000110101000110,
16'b1000110110111001,
16'b1000111000101101,
16'b1000111010100011,
16'b1000111100011011,
16'b1000111110010100,
16'b1001000000001111,
16'b1001000010001100,
16'b1001000100001011,
16'b1001000110001100,
16'b1001001000001110,
16'b1001001010010010,
16'b1001001100011000,
16'b1001001110011111,
16'b1001010000101000,
16'b1001010010110011,
16'b1001010100111111,
16'b1001010111001101,
16'b1001011001011101,
16'b1001011011101110,
16'b1001011110000001,
16'b1001100000010110,
16'b1001100010101100,
16'b1001100101000100,
16'b1001100111011110,
16'b1001101001111001,
16'b1001101100010110,
16'b1001101110110100,
16'b1001110001010100,
16'b1001110011110101,
16'b1001110110011000,
16'b1001111000111101,
16'b1001111011100011,
16'b1001111110001010,
16'b1010000000110011,
16'b1010000011011110,
16'b1010000110001010,
16'b1010001000110111,
16'b1010001011100110,
16'b1010001110010110,
16'b1010010001001000,
16'b1010010011111100,
16'b1010010110110000,
16'b1010011001100110,
16'b1010011100011110,
16'b1010011111010111,
16'b1010100010010001,
16'b1010100101001101,
16'b1010101000001010,
16'b1010101011001000,
16'b1010101110001000,
16'b1010110001001001,
16'b1010110100001011,
16'b1010110111001111,
16'b1010111010010100,
16'b1010111101011010,
16'b1011000000100001,
16'b1011000011101010,
16'b1011000110110100,
16'b1011001001111111,
16'b1011001101001011,
16'b1011010000011001,
16'b1011010011101000,
16'b1011010110111000,
16'b1011011010001001,
16'b1011011101011011,
16'b1011100000101110,
16'b1011100100000011,
16'b1011100111011000,
16'b1011101010101111,
16'b1011101110000111,
16'b1011110001011111,
16'b1011110100111001,
16'b1011111000010100,
16'b1011111011110000,
16'b1011111111001101,
16'b1100000010101011,
16'b1100000110001010,
16'b1100001001101010,
16'b1100001101001011,
16'b1100010000101101,
16'b1100010100010000,
16'b1100010111110011,
16'b1100011011011000,
16'b1100011110111101,
16'b1100100010100100,
16'b1100100110001011,
16'b1100101001110011,
16'b1100101101011100,
16'b1100110001000110,
16'b1100110100110000,
16'b1100111000011100,
16'b1100111100001000,
16'b1100111111110101,
16'b1101000011100010,
16'b1101000111010001,
16'b1101001011000000,
16'b1101001110110000,
16'b1101010010100000,
16'b1101010110010010,
16'b1101011010000011,
16'b1101011101110110,
16'b1101100001101001,
16'b1101100101011101,
16'b1101101001010001,
16'b1101101101000110,
16'b1101110000111100,
16'b1101110100110010,
16'b1101111000101000,
16'b1101111100011111,
16'b1110000000010111,
16'b1110000100001111,
16'b1110001000001000,
16'b1110001100000001,
16'b1110001111111011,
16'b1110010011110101,
16'b1110010111101111,
16'b1110011011101010,
16'b1110011111100101,
16'b1110100011100001,
16'b1110100111011101,
16'b1110101011011001,
16'b1110101111010110,
16'b1110110011010011,
16'b1110110111010000,
16'b1110111011001101,
16'b1110111111001011,
16'b1111000011001001,
16'b1111000111001000,
16'b1111001011000110,
16'b1111001111000101,
16'b1111010011000100,
16'b1111010111000011,
16'b1111011011000010,
16'b1111011111000010,
16'b1111100011000001,
16'b1111100111000001,
16'b1111101011000000,
16'b1111101111000000,
16'b1111110011000000,
16'b1111110111000000,
16'b1111111011000000,
16'b1111111111000000,
16'b0000000011000000,
16'b0000000111000000,
16'b0000001011000000,
16'b0000001111000000,
16'b0000010011000000,
16'b0000010111000000,
16'b0000011010111111,
16'b0000011110111111,
16'b0000100010111110,
16'b0000100110111110,
16'b0000101010111101,
16'b0000101110111100,
16'b0000110010111011,
16'b0000110110111001,
16'b0000111010111000,
16'b0000111110110110,
16'b0001000010110100,
16'b0001000110110010,
16'b0001001010101111,
16'b0001001110101100,
16'b0001010010101001,
16'b0001010110100101,
16'b0001011010100001,
16'b0001011110011101,
16'b0001100010011001,
16'b0001100110010100,
16'b0001101010001110,
16'b0001101110001001,
16'b0001110010000010,
16'b0001110101111100,
16'b0001111001110101,
16'b0001111101101101,
16'b0010000001100101,
16'b0010000101011100,
16'b0010001001010011,
16'b0010001101001010,
16'b0010010000111111,
16'b0010010100110101,
16'b0010011000101001,
16'b0010011100011101,
16'b0010100000010001,
16'b0010100100000100,
16'b0010100111110110,
16'b0010101011100111,
16'b0010101111011000,
16'b0010110011001000,
16'b0010110110111000,
16'b0010111010100110,
16'b0010111110010101,
16'b0011000010000010,
16'b0011000101101110,
16'b0011001001011010,
16'b0011001101000101,
16'b0011010000101111,
16'b0011010100011001,
16'b0011011000000001,
16'b0011011011101001,
16'b0011011111010000,
16'b0011100010110101,
16'b0011100110011011,
16'b0011101001111111,
16'b0011101101100010,
16'b0011110001000100,
16'b0011110100100110,
16'b0011111000000110,
16'b0011111011100110,
16'b0011111111000100,
16'b0100000010100001,
16'b0100000101111110,
16'b0100001001011001,
16'b0100001100110100,
16'b0100010000001101,
16'b0100010011100101,
16'b0100010110111101,
16'b0100011010010011,
16'b0100011101101000,
16'b0100100000111100,
16'b0100100100001110,
16'b0100100111100000,
16'b0100101010110001,
16'b0100101110000000,
16'b0100110001001110,
16'b0100110100011011,
16'b0100110111100111,
16'b0100111010110001,
16'b0100111101111010,
16'b0101000001000010,
16'b0101000100001001,
16'b0101000111001111,
16'b0101001010010011,
16'b0101001101010110,
16'b0101010000011000,
16'b0101010011011000,
16'b0101010110010111,
16'b0101011001010101,
16'b0101011100010001,
16'b0101011111001100,
16'b0101100010000110,
16'b0101100100111110,
16'b0101100111110101,
16'b0101101010101010,
16'b0101101101011110,
16'b0101110000010001,
16'b0101110011000010,
16'b0101110101110001,
16'b0101111000100000,
16'b0101111011001100,
16'b0101111101111000,
16'b0110000000100001,
16'b0110000011001010,
16'b0110000101110000,
16'b0110001000010110,
16'b0110001010111001,
16'b0110001101011100,
16'b0110001111111100,
16'b0110010010011011,
16'b0110010100111001,
16'b0110010111010101,
16'b0110011001101111,
16'b0110011100001000,
16'b0110011110011111,
16'b0110100000110100,
16'b0110100011001000,
16'b0110100101011010,
16'b0110100111101011,
16'b0110101001111010,
16'b0110101100000111,
16'b0110101110010011,
16'b0110110000011100,
16'b0110110010100101,
16'b0110110100101011,
16'b0110110110110000,
16'b0110111000110011,
16'b0110111010110100,
16'b0110111100110100,
16'b0110111110110010,
16'b0111000000101110,
16'b0111000010101000,
16'b0111000100100001,
16'b0111000110011000,
16'b0111001000001101,
16'b0111001010000000,
16'b0111001011110010,
16'b0111001101100010,
16'b0111001111010000,
16'b0111010000111100,
16'b0111010010100110,
16'b0111010100001110,
16'b0111010101110101,
16'b0111010111011010,
16'b0111011000111101,
16'b0111011010011110,
16'b0111011011111101,
16'b0111011101011011,
16'b0111011110110110,
16'b0111100000010000,
16'b0111100001101000,
16'b0111100010111110,
16'b0111100100010010,
16'b0111100101100100,
16'b0111100110110100,
16'b0111101000000010,
16'b0111101001001111,
16'b0111101010011001,
16'b0111101011100010,
16'b0111101100101001,
16'b0111101101101101,
16'b0111101110110000,
16'b0111101111110001,
16'b0111110000110000,
16'b0111110001101101,
16'b0111110010101000,
16'b0111110011100001,
16'b0111110100011001,
16'b0111110101001110,
16'b0111110110000001,
16'b0111110110110010,
16'b0111110111100010,
16'b0111111000001111,
16'b0111111000111010,
16'b0111111001100100,
16'b0111111010001011,
16'b0111111010110001,
16'b0111111011010100,
16'b0111111011110110,
16'b0111111100010101,
16'b0111111100110011,
16'b0111111101001111,
16'b0111111101101000,
16'b0111111110000000,
16'b0111111110010101,
16'b0111111110101001,
16'b0111111110111010,
16'b0111111111001010,
16'b0111111111011000,
16'b0111111111100011,
16'b0111111111101101,
16'b0111111111110101,
16'b0111111111111010,
16'b0111111111111110,
16'b0111111111111111,
16'b0111111111111111,
16'b0111111111111101,
16'b0111111111111000,
16'b0111111111110010,
16'b0111111111101010,
16'b0111111111011111,
16'b0111111111010011,
16'b0111111111000100,
16'b0111111110110100,
16'b0111111110100010,
16'b0111111110001101,
16'b0111111101110111,
16'b0111111101011111,
16'b0111111101000100,
16'b0111111100101000,
16'b0111111100001010,
16'b0111111011101001,
16'b0111111011000111
};

assign out = ROM[theta];

endmodule